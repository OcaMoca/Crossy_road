
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity ram is
	generic
	(
		DATA_WIDTH : natural := 32;		    -- 4 byte one line of memory
		ADDR_WIDTH : natural := 13			    -- 24576 bytes size of memory
	);

	port(
		i_clk    : in  std_logic;
		i_r_addr : in  std_logic_vector(ADDR_WIDTH-1 downto 0);
		i_data   : in  std_logic_vector(DATA_WIDTH-1 downto 0);
		i_we     : in  std_logic;
		i_w_addr : in  std_logic_vector(ADDR_WIDTH-1 downto 0);
		o_data   : out std_logic_vector(DATA_WIDTH-1 downto 0)
	);
end entity ram;

architecture arch of ram is

	type ram_t is array (0 to 2**ADDR_WIDTH-1) of std_logic_vector(DATA_WIDTH-1 downto 0);


-- GENERATED BY BC_MEM_PACKER

-- DATE: Thu May 18 16:01:02 2017

	signal mem : ram_t := (

--			***** COLOR PALLETE *****


--kirby colors
        0 => x"00000000",
        1=> x"00ea8bff",
        2 => x"00e98afe",
        3 => x"003d3d40",
        4 => x"00811699",
        5 => x"00ea8aff",
        6 => x"000303d5",
--mapa colors
	7=> x"00353b39",
	8=> x"000cac83",
	9=> x"00ffffff",
	10=> x"009b6f2e",
	11=> x"00000000",
	12=> x"0019704d",
	13=> x"00010101",
	14=> x"001b714d",
	15=> x"001b714e",
	16=> x"001c714e",
	17=> x"001a6e4f",
	
--deblo
	 18 =>x"00000000
         19 =>x"0008072c
         
--red_car
          
                20=> x"00000000",
                21=> x"00000001",
                22=> x"00000002",
                23=> x"00010104",
                24=> x"0007072c",
                25=> x"0002020c",
                26=> x"00010102",
                27=> x"00020001",
                28=> x"000000fe",
                29=> x"0008072c",
                30=> x"00b19357",
                31=> x"000800fe",
                32=> x"0000dcd6",
                33=> x"0012082c",
                34=> x"0019092c",
                35=> x"0016092c",
                36=> x"001d01fb",
                37=> x"00000003",
                38=> x"00010001",
                
--blue_car
                
        39=> x"00000000",
        40=> x"00000001",
        41=> x"00000002",
        42=> x"0008072c",
        43=> x"00070102",
        44=> x"00020102",
        45=> x"00010002",
        46=> x"00ab1c2b",
        47=> x"00b09256",
        48=> x"0000dcd6",
        49=> x"000e082c",
        50=> x"00020101",
        51=> x"00010000",
        52=> x"00060102",
        53=> x"00010102",     
                


            --  ADDED SPRITES HERE
          --  SPRITE
		64 => x"0202020F",
		65 => x"3C020202",
		66 => x"02020202",
		67 => x"02020202",
		68 => x"02020F0F",
		69 => x"3C3C0202",
		70 => x"02020202",
		71 => x"02020202",
		72 => x"020F0F0F",
		73 => x"3C3C3C02",
		74 => x"02020202",
		75 => x"02020202",
		76 => x"0F3C0F3C",
		77 => x"023C023C",
		78 => x"02020202",
		79 => x"02020202",
		80 => x"0F0F3C3C",
		81 => x"3C023C3C",
		82 => x"02020202",
		83 => x"02020202",
		84 => x"0F0F3C3C",
		85 => x"3C023C3C",
		86 => x"02020202",
		87 => x"02020202",
		88 => x"0F0F3C3C",
		89 => x"3C023C3C",
		90 => x"02020202",
		91 => x"02020202",
		92 => x"0F0F3C3C",
		93 => x"3C023C3C",
		94 => x"02020202",
		95 => x"02020202",
		96 => x"0F0F3C3C",
		97 => x"3C023C3C",
		98 => x"02020202",
		99 => x"02020202",
		100 => x"0F0F3C3C",
		101 => x"3C023C3C",
		102 => x"02020202",
		103 => x"02020202",
		104 => x"0F0F3C3C",
		105 => x"3C023C3C",
		106 => x"02020202",
		107 => x"02020202",
		108 => x"0F3C0F3C",
		109 => x"3C023C3C",
		110 => x"02020202",
		111 => x"02020202",
		112 => x"3C3C3C0F",
		113 => x"023C023C",
		114 => x"02020202",
		115 => x"02020202",
		116 => x"023C3C3C",
		117 => x"3C3C3C02",
		118 => x"02020202",
		119 => x"02020202",
		120 => x"02023C3C",
		121 => x"3C3C0202",
		122 => x"02020202",
		123 => x"02020202",
		124 => x"0202023C",
		125 => x"3C020202",
		126 => x"02020202",
		127 => x"02020202",

          -- BOMB SPRITE
		128 => x"02020202",
		129 => x"020F0202",
		130 => x"02020202",
		131 => x"02020202",
		132 => x"02020202",
		133 => x"020F0202",
		134 => x"02020202",
		135 => x"02020202",
		136 => x"02020202",
		137 => x"02020F02",
		138 => x"02020202",
		139 => x"02020202",
		140 => x"02020202",
		141 => x"0202020F",
		142 => x"02020202",
		143 => x"02020202",
		144 => x"02020202",
		145 => x"0202020F",
		146 => x"02020202",
		147 => x"02020202",
		148 => x"02020202",
		149 => x"02020F02",
		150 => x"02020202",
		151 => x"02020202",
		152 => x"02020D0D",
		153 => x"0D0D0202",
		154 => x"02020202",
		155 => x"02020202",
		156 => x"020D2E2E",
		157 => x"0D0D0D02",
		158 => x"02020202",
		159 => x"02020202",
		160 => x"0D2E0F2E",
		161 => x"0D0D0D0D",
		162 => x"02020202",
		163 => x"02020202",
		164 => x"0D2E2E0D",
		165 => x"0D0D0D0D",
		166 => x"02020202",
		167 => x"02020202",
		168 => x"0D0D0D0D",
		169 => x"0D0D0D0D",
		170 => x"02020202",
		171 => x"02020202",
		172 => x"0D0D0D0D",
		173 => x"0D0D0D0D",
		174 => x"02020202",
		175 => x"02020202",
		176 => x"020D0D0D",
		177 => x"0D0D0D02",
		178 => x"02020202",
		179 => x"02020202",
		180 => x"02020D0D",
		181 => x"0D0D0202",
		182 => x"02020202",
		183 => x"02020202",
		184 => x"02020202",
		185 => x"02020202",
		186 => x"02020202",
		187 => x"02020202",
		188 => x"02020202",
		189 => x"02020202",
		190 => x"02020202",
		191 => x"02020202",

--			***** 16x16 IMAGES *****
--			OVERWORLD SPRITES
        
        --kirby sprites        
               
                --  sprite 0
        255 => x"08080808",		-- colors: 8, 8, 8, 8
        256 => x"08080808",		-- colors: 8, 8, 8, 8
        257 => x"08080808",		-- colors: 8, 8, 8, 8
        258 => x"08080808",		-- colors: 8, 8, 8, 8
        259 => x"08080808",		-- colors: 8, 8, 8, 8
        260 => x"08080808",		-- colors: 8, 8, 8, 8
        261 => x"08080808",		-- colors: 8, 8, 8, 8
        262 => x"08080808",		-- colors: 8, 8, 8, 8
        263 => x"08080808",		-- colors: 8, 8, 8, 8
        264 => x"08080808",		-- colors: 8, 8, 8, 8
        265 => x"08080808",		-- colors: 8, 8, 8, 8
        266 => x"08080808",		-- colors: 8, 8, 8, 8
        267 => x"08080808",		-- colors: 8, 8, 8, 8
        268 => x"08080808",		-- colors: 8, 8, 8, 8
        269 => x"08080808",		-- colors: 8, 8, 8, 8
        270 => x"08080808",		-- colors: 8, 8, 8, 8
        271 => x"08080808",		-- colors: 8, 8, 8, 8
        272 => x"08080808",		-- colors: 8, 8, 8, 8
        273 => x"08080808",		-- colors: 8, 8, 8, 8
        274 => x"08080808",		-- colors: 8, 8, 8, 8
        275 => x"08080808",		-- colors: 8, 8, 8, 8
        276 => x"08080808",		-- colors: 8, 8, 8, 8
        277 => x"08080808",		-- colors: 8, 8, 8, 8
        278 => x"08080808",		-- colors: 8, 8, 8, 8
        279 => x"08080808",		-- colors: 8, 8, 8, 8
        280 => x"08080808",		-- colors: 8, 8, 8, 8
        281 => x"08080808",		-- colors: 8, 8, 8, 8
        282 => x"08080808",		-- colors: 8, 8, 8, 8
        283 => x"08080808",		-- colors: 8, 8, 8, 8
        284 => x"08080909",		-- colors: 8, 8, 9, 9
        285 => x"090A0808",		-- colors: 9, 10, 8, 8
        286 => x"08080808",		-- colors: 8, 8, 8, 8
        287 => x"08080808",		-- colors: 8, 8, 8, 8
        288 => x"08090909",		-- colors: 8, 9, 9, 9
        289 => x"09090908",		-- colors: 9, 9, 9, 8
        290 => x"08080808",		-- colors: 8, 8, 8, 8
        291 => x"08080808",		-- colors: 8, 8, 8, 8
        292 => x"09090B09",		-- colors: 9, 9, 11, 9
        293 => x"090B0909",		-- colors: 9, 11, 9, 9
        294 => x"08080808",		-- colors: 8, 8, 8, 8
        295 => x"08080809",		-- colors: 8, 8, 8, 9
        296 => x"09090B09",		-- colors: 9, 9, 11, 9
        297 => x"090B0909",		-- colors: 9, 11, 9, 9
        298 => x"09080808",		-- colors: 9, 8, 8, 8
        299 => x"08080809",		-- colors: 8, 8, 8, 9
        300 => x"090C0909",		-- colors: 9, 12, 9, 9
        301 => x"09090C09",		-- colors: 9, 9, 12, 9
        302 => x"09080808",		-- colors: 9, 8, 8, 8
        303 => x"08080808",		-- colors: 8, 8, 8, 8
        304 => x"0D090909",		-- colors: 13, 9, 9, 9
        305 => x"09090909",		-- colors: 9, 9, 9, 9
        306 => x"08080808",		-- colors: 8, 8, 8, 8
        307 => x"08080808",		-- colors: 8, 8, 8, 8
        308 => x"08090909",		-- colors: 8, 9, 9, 9
        309 => x"09090908",		-- colors: 9, 9, 9, 8
        310 => x"08080808",		-- colors: 8, 8, 8, 8
        311 => x"08080808",		-- colors: 8, 8, 8, 8
        312 => x"08080909",		-- colors: 8, 8, 9, 9
        313 => x"09090808",		-- colors: 9, 9, 8, 8
        314 => x"08080808",		-- colors: 8, 8, 8, 8
        315 => x"08080808",		-- colors: 8, 8, 8, 8
        316 => x"080E0E08",		-- colors: 8, 14, 14, 8
        317 => x"080E0E08",		-- colors: 8, 14, 14, 8
        318 => x"08080808",		-- colors: 8, 8, 8, 8
        
        --deblo sprite
        
                --  sprite 0
        319 => x"2E2E2E2E",		-- colors: 46, 46, 46, 46
        320 => x"2E2E2E2E",		-- colors: 46, 46, 46, 46
        321 => x"2E2E2E2E",		-- colors: 46, 46, 46, 46
        322 => x"2E2E2E2E",		-- colors: 46, 46, 46, 46
        323 => x"2E2E2E2E",		-- colors: 46, 46, 46, 46
        324 => x"2E2E2E2E",		-- colors: 46, 46, 46, 46
        325 => x"2E2E2E2E",		-- colors: 46, 46, 46, 46
        326 => x"2E2E2E2E",		-- colors: 46, 46, 46, 46
        327 => x"2E2E2E2E",		-- colors: 46, 46, 46, 46
        328 => x"2E2E2E2E",		-- colors: 46, 46, 46, 46
        329 => x"2E2E2E2E",		-- colors: 46, 46, 46, 46
        330 => x"2E2E2E2E",		-- colors: 46, 46, 46, 46
        331 => x"2E2E2E2E",		-- colors: 46, 46, 46, 46
        332 => x"2E2E2E2E",		-- colors: 46, 46, 46, 46
        333 => x"2E2E2E2E",		-- colors: 46, 46, 46, 46
        334 => x"2E2E2E2E",		-- colors: 46, 46, 46, 46
        335 => x"2E2E2E2E",		-- colors: 46, 46, 46, 46
        336 => x"2E2E2E2E",		-- colors: 46, 46, 46, 46
        337 => x"2E2E2E2E",		-- colors: 46, 46, 46, 46
        338 => x"2E2E2E2E",		-- colors: 46, 46, 46, 46
        339 => x"2E2E2E2E",		-- colors: 46, 46, 46, 46
        340 => x"2E2E2E2E",		-- colors: 46, 46, 46, 46
        341 => x"2E2E2E2E",		-- colors: 46, 46, 46, 46
        342 => x"2E2E2E2E",		-- colors: 46, 46, 46, 46
        343 => x"2E2E2E2E",		-- colors: 46, 46, 46, 46
        344 => x"2E2E2E2E",		-- colors: 46, 46, 46, 46
        345 => x"2E2E2E2E",		-- colors: 46, 46, 46, 46
        346 => x"2E2E2E2E",		-- colors: 46, 46, 46, 46
        347 => x"2F2F2F2F",		-- colors: 47, 47, 47, 47
        348 => x"2F2F2F2F",		-- colors: 47, 47, 47, 47
        349 => x"2F2F2F2F",		-- colors: 47, 47, 47, 47
        350 => x"2F2F2F2F",		-- colors: 47, 47, 47, 47
        351 => x"2F2F2F2F",		-- colors: 47, 47, 47, 47
        352 => x"2F2F2F2F",		-- colors: 47, 47, 47, 47
        353 => x"2F2F2F2F",		-- colors: 47, 47, 47, 47
        354 => x"2F2F2F2F",		-- colors: 47, 47, 47, 47
        355 => x"2F2F2F2F",		-- colors: 47, 47, 47, 47
        356 => x"2F2F2F2F",		-- colors: 47, 47, 47, 47
        357 => x"2F2F2F2F",		-- colors: 47, 47, 47, 47
        358 => x"2F2F2F2F",		-- colors: 47, 47, 47, 47
        359 => x"2F2F2F2F",		-- colors: 47, 47, 47, 47
        360 => x"2F2F2F2F",		-- colors: 47, 47, 47, 47
        361 => x"2F2F2F2F",		-- colors: 47, 47, 47, 47
        362 => x"2F2F2F2F",		-- colors: 47, 47, 47, 47
        363 => x"2F2F2F2F",		-- colors: 47, 47, 47, 47
        364 => x"2F2F2F2F",		-- colors: 47, 47, 47, 47
        365 => x"2F2F2F2F",		-- colors: 47, 47, 47, 47
        366 => x"2F2F2F2F",		-- colors: 47, 47, 47, 47
        367 => x"2F2F2F2F",		-- colors: 47, 47, 47, 47
        368 => x"2F2F2F2F",		-- colors: 47, 47, 47, 47
        369 => x"2F2F2F2F",		-- colors: 47, 47, 47, 47
        370 => x"2F2F2F2F",		-- colors: 47, 47, 47, 47
        371 => x"2F2F2F2F",		-- colors: 47, 47, 47, 47
        372 => x"2F2F2F2F",		-- colors: 47, 47, 47, 47
        373 => x"2F2F2F2F",		-- colors: 47, 47, 47, 47
        374 => x"2F2F2F2F",		-- colors: 47, 47, 47, 47
        375 => x"2F2F2F2F",		-- colors: 47, 47, 47, 47
        376 => x"2F2F2F2F",		-- colors: 47, 47, 47, 47
        377 => x"2F2F2F2F",		-- colors: 47, 47, 47, 47
        378 => x"2F2F2F2F",		-- colors: 47, 47, 47, 47
        379 => x"2F2F2F2F",		-- colors: 47, 47, 47, 47
        380 => x"2F2F2F2F",		-- colors: 47, 47, 47, 47
        381 => x"2F2F2F2F",		-- colors: 47, 47, 47, 47
        382 => x"2F2F2F2F",		-- colors: 47, 47, 47, 47

                --  sprite 1
        383 => x"2E2E2E2E",		-- colors: 46, 46, 46, 46
        384 => x"2E2E2E2E",		-- colors: 46, 46, 46, 46
        385 => x"2E2E2E2E",		-- colors: 46, 46, 46, 46
        386 => x"2E2E2E2E",		-- colors: 46, 46, 46, 46
        387 => x"2E2E2E2E",		-- colors: 46, 46, 46, 46
        388 => x"2E2E2E2E",		-- colors: 46, 46, 46, 46
        389 => x"2E2E2E2E",		-- colors: 46, 46, 46, 46
        390 => x"2E2E2E2E",		-- colors: 46, 46, 46, 46
        391 => x"2E2E2E2E",		-- colors: 46, 46, 46, 46
        392 => x"2E2E2E2E",		-- colors: 46, 46, 46, 46
        393 => x"2E2E2E2E",		-- colors: 46, 46, 46, 46
        394 => x"2E2E2E2E",		-- colors: 46, 46, 46, 46
        395 => x"2E2E2E2E",		-- colors: 46, 46, 46, 46
        396 => x"2E2E2E2E",		-- colors: 46, 46, 46, 46
        397 => x"2E2E2E2E",		-- colors: 46, 46, 46, 46
        398 => x"2E2E2E2E",		-- colors: 46, 46, 46, 46
        399 => x"2E2E2E2E",		-- colors: 46, 46, 46, 46
        400 => x"2E2E2E2E",		-- colors: 46, 46, 46, 46
        401 => x"2E2E2E2E",		-- colors: 46, 46, 46, 46
        402 => x"2E2E2E2E",		-- colors: 46, 46, 46, 46
        403 => x"2E2E2E2E",		-- colors: 46, 46, 46, 46
        404 => x"2E2E2E2E",		-- colors: 46, 46, 46, 46
        405 => x"2E2E2E2E",		-- colors: 46, 46, 46, 46
        406 => x"2E2E2E2E",		-- colors: 46, 46, 46, 46
        407 => x"2E2E2E2E",		-- colors: 46, 46, 46, 46
        408 => x"2E2E2E2E",		-- colors: 46, 46, 46, 46
        409 => x"2E2E2E2E",		-- colors: 46, 46, 46, 46
        410 => x"2E2E2E2E",		-- colors: 46, 46, 46, 46
        411 => x"2F2F2F2F",		-- colors: 47, 47, 47, 47
        412 => x"2F2F2F2F",		-- colors: 47, 47, 47, 47
        413 => x"2F2F2F2F",		-- colors: 47, 47, 47, 47
        414 => x"2F2F2F2F",		-- colors: 47, 47, 47, 47
        415 => x"2F2F2F2F",		-- colors: 47, 47, 47, 47
        416 => x"2F2F2F2F",		-- colors: 47, 47, 47, 47
        417 => x"2F2F2F2F",		-- colors: 47, 47, 47, 47
        418 => x"2F2F2F2F",		-- colors: 47, 47, 47, 47
        419 => x"2F2F2F2F",		-- colors: 47, 47, 47, 47
        420 => x"2F2F2F2F",		-- colors: 47, 47, 47, 47
        421 => x"2F2F2F2F",		-- colors: 47, 47, 47, 47
        422 => x"2F2F2F2F",		-- colors: 47, 47, 47, 47
        423 => x"2F2F2F2F",		-- colors: 47, 47, 47, 47
        424 => x"2F2F2F2F",		-- colors: 47, 47, 47, 47
        425 => x"2F2F2F2F",		-- colors: 47, 47, 47, 47
        426 => x"2F2F2F2F",		-- colors: 47, 47, 47, 47
        427 => x"2F2F2F2F",		-- colors: 47, 47, 47, 47
        428 => x"2F2F2F2F",		-- colors: 47, 47, 47, 47
        429 => x"2F2F2F2F",		-- colors: 47, 47, 47, 47
        430 => x"2F2F2F2F",		-- colors: 47, 47, 47, 47
        431 => x"2F2F2F2F",		-- colors: 47, 47, 47, 47
        432 => x"2F2F2F2F",		-- colors: 47, 47, 47, 47
        433 => x"2F2F2F2F",		-- colors: 47, 47, 47, 47
        434 => x"2F2F2F2F",		-- colors: 47, 47, 47, 47
        435 => x"2F2F2F2F",		-- colors: 47, 47, 47, 47
        436 => x"2F2F2F2F",		-- colors: 47, 47, 47, 47
        437 => x"2F2F2F2F",		-- colors: 47, 47, 47, 47
        438 => x"2F2F2F2F",		-- colors: 47, 47, 47, 47
        439 => x"2F2F2F2F",		-- colors: 47, 47, 47, 47
        440 => x"2F2F2F2F",		-- colors: 47, 47, 47, 47
        441 => x"2F2F2F2F",		-- colors: 47, 47, 47, 47
        442 => x"2F2F2F2F",		-- colors: 47, 47, 47, 47
        443 => x"2F2F2F2F",		-- colors: 47, 47, 47, 47
        444 => x"2F2F2F2F",		-- colors: 47, 47, 47, 47
        445 => x"2F2F2F2F",		-- colors: 47, 47, 47, 47
        446 => x"2F2F2F2F",		-- colors: 47, 47, 47, 47

        
--red_car sprite



                --  sprite 0
        447 => x"14141414",		-- colors: 20, 20, 20, 20
        448 => x"14141516",		-- colors: 20, 20, 21, 22
        449 => x"16161515",		-- colors: 22, 22, 21, 21
        450 => x"15141414",		-- colors: 21, 20, 20, 20
        451 => x"14141414",		-- colors: 20, 20, 20, 20
        452 => x"14171818",		-- colors: 20, 23, 24, 24
        453 => x"18181815",		-- colors: 24, 24, 24, 21
        454 => x"15151515",		-- colors: 21, 21, 21, 21
        455 => x"14141415",		-- colors: 20, 20, 20, 21
        456 => x"16191818",		-- colors: 22, 25, 24, 24
        457 => x"18181818",		-- colors: 24, 24, 24, 24
        458 => x"151A151B",		-- colors: 21, 26, 21, 27
        459 => x"14151818",		-- colors: 20, 21, 24, 24
        460 => x"18181818",		-- colors: 24, 24, 24, 24
        461 => x"1C1C1C1C",		-- colors: 28, 28, 28, 28
        462 => x"1D1D1C1C",		-- colors: 29, 29, 28, 28
        463 => x"1618181C",		-- colors: 22, 24, 24, 28
        464 => x"1C1C1818",		-- colors: 28, 28, 24, 24
        465 => x"1C1C1C1C",		-- colors: 28, 28, 28, 28
        466 => x"1D1D1C1C",		-- colors: 29, 29, 28, 28
        467 => x"18181F1C",		-- colors: 24, 24, 31, 28
        468 => x"1C1C1818",		-- colors: 28, 28, 24, 24
        469 => x"1D1D1D1D",		-- colors: 29, 29, 29, 29
        470 => x"1D1D1D1D",		-- colors: 29, 29, 29, 29
        471 => x"18181C1C",		-- colors: 24, 24, 28, 28
        472 => x"1C1C1818",		-- colors: 28, 28, 24, 24
        473 => x"1C1C1C1C",		-- colors: 28, 28, 28, 28
        474 => x"1C1C1C1C",		-- colors: 28, 28, 28, 28
        475 => x"18181C1C",		-- colors: 24, 24, 28, 28
        476 => x"1C1C1818",		-- colors: 28, 28, 24, 24
        477 => x"1C1C1C1C",		-- colors: 28, 28, 28, 28
        478 => x"1C1C1C1D",		-- colors: 28, 28, 28, 29
        479 => x"18181C1C",		-- colors: 24, 24, 28, 28
        480 => x"1C1C1818",		-- colors: 28, 28, 24, 24
        481 => x"1C1C1C1C",		-- colors: 28, 28, 28, 28
        482 => x"1C1C1C1C",		-- colors: 28, 28, 28, 28
        483 => x"18181C1C",		-- colors: 24, 24, 28, 28
        484 => x"1C1C1818",		-- colors: 28, 28, 24, 24
        485 => x"21222223",		-- colors: 33, 34, 34, 35
        486 => x"1D1D1D1D",		-- colors: 29, 29, 29, 29
        487 => x"1518181C",		-- colors: 21, 24, 24, 28
        488 => x"1C1C1818",		-- colors: 28, 28, 24, 24
        489 => x"1C1C1C1C",		-- colors: 28, 28, 28, 28
        490 => x"1D1D1C1C",		-- colors: 29, 29, 28, 28
        491 => x"15251818",		-- colors: 21, 37, 24, 24
        492 => x"18181818",		-- colors: 24, 24, 24, 24
        493 => x"1C1C1C1C",		-- colors: 28, 28, 28, 28
        494 => x"1D1D1C1C",		-- colors: 29, 29, 28, 28
        495 => x"15151515",		-- colors: 21, 21, 21, 21
        496 => x"16151818",		-- colors: 22, 21, 24, 24
        497 => x"18181818",		-- colors: 24, 24, 24, 24
        498 => x"14152626",		-- colors: 20, 21, 38, 38
        499 => x"14141515",		-- colors: 20, 20, 21, 21
        500 => x"14151818",		-- colors: 20, 21, 24, 24
        501 => x"18181814",		-- colors: 24, 24, 24, 20
        502 => x"15141414",		-- colors: 21, 20, 20, 20
        503 => x"14141414",		-- colors: 20, 20, 20, 20
        504 => x"14141415",		-- colors: 20, 20, 20, 21
        505 => x"16161514",		-- colors: 22, 22, 21, 20
        506 => x"14141414",		-- colors: 20, 20, 20, 20
        507 => x"14141414",		-- colors: 20, 20, 20, 20
        508 => x"14141414",		-- colors: 20, 20, 20, 20
        509 => x"14141414",		-- colors: 20, 20, 20, 20
        510 => x"14141414",		-- colors: 20, 20, 20, 20

                --  sprite 1
        511 => x"14141414",		-- colors: 20, 20, 20, 20
        512 => x"14141414",		-- colors: 20, 20, 20, 20
        513 => x"14141414",		-- colors: 20, 20, 20, 20
        514 => x"14141414",		-- colors: 20, 20, 20, 20
        515 => x"14151818",		-- colors: 20, 21, 24, 24
        516 => x"18181818",		-- colors: 24, 24, 24, 24
        517 => x"18151514",		-- colors: 24, 21, 21, 20
        518 => x"14141414",		-- colors: 20, 20, 20, 20
        519 => x"18181818",		-- colors: 24, 24, 24, 24
        520 => x"18181818",		-- colors: 24, 24, 24, 24
        521 => x"18181515",		-- colors: 24, 24, 21, 21
        522 => x"15141414",		-- colors: 21, 20, 20, 20
        523 => x"18181E1E",		-- colors: 24, 24, 30, 30
        524 => x"1C1C1C1C",		-- colors: 28, 28, 28, 28
        525 => x"1C1C1818",		-- colors: 28, 28, 24, 24
        526 => x"15161514",		-- colors: 21, 22, 21, 20
        527 => x"18181E1E",		-- colors: 24, 24, 30, 30
        528 => x"1E1E1C1C",		-- colors: 30, 30, 28, 28
        529 => x"1C1C1C1C",		-- colors: 28, 28, 28, 28
        530 => x"18181515",		-- colors: 24, 24, 21, 21
        531 => x"18181E1E",		-- colors: 24, 24, 30, 30
        532 => x"1E1E1E1E",		-- colors: 30, 30, 30, 30
        533 => x"1C1C1C1C",		-- colors: 28, 28, 28, 28
        534 => x"1C1C2020",		-- colors: 28, 28, 32, 32
        535 => x"18181E1E",		-- colors: 24, 24, 30, 30
        536 => x"1E1E1E1E",		-- colors: 30, 30, 30, 30
        537 => x"1E1C1C1C",		-- colors: 30, 28, 28, 28
        538 => x"1C1C1818",		-- colors: 28, 28, 24, 24
        539 => x"18181E1E",		-- colors: 24, 24, 30, 30
        540 => x"1E1E1E1E",		-- colors: 30, 30, 30, 30
        541 => x"1E1C1C1C",		-- colors: 30, 28, 28, 28
        542 => x"1C1C1818",		-- colors: 28, 28, 24, 24
        543 => x"18181E1E",		-- colors: 24, 24, 30, 30
        544 => x"1E1E1E1E",		-- colors: 30, 30, 30, 30
        545 => x"1E1C1C1C",		-- colors: 30, 28, 28, 28
        546 => x"1C1C1818",		-- colors: 28, 28, 24, 24
        547 => x"18181E1E",		-- colors: 24, 24, 30, 30
        548 => x"1E1E1E1E",		-- colors: 30, 30, 30, 30
        549 => x"1C1C1C1C",		-- colors: 28, 28, 28, 28
        550 => x"1C1C2020",		-- colors: 28, 28, 32, 32
        551 => x"18181E1E",		-- colors: 24, 24, 30, 30
        552 => x"1E1E241C",		-- colors: 30, 30, 36, 28
        553 => x"1C1C1C1C",		-- colors: 28, 28, 28, 28
        554 => x"18181515",		-- colors: 24, 24, 21, 21
        555 => x"18181E1E",		-- colors: 24, 24, 30, 30
        556 => x"1C1C1C1C",		-- colors: 28, 28, 28, 28
        557 => x"1C1C1818",		-- colors: 28, 28, 24, 24
        558 => x"15161515",		-- colors: 21, 22, 21, 21
        559 => x"18181818",		-- colors: 24, 24, 24, 24
        560 => x"18181818",		-- colors: 24, 24, 24, 24
        561 => x"18181515",		-- colors: 24, 24, 21, 21
        562 => x"16141414",		-- colors: 22, 20, 20, 20
        563 => x"14151818",		-- colors: 20, 21, 24, 24
        564 => x"18181818",		-- colors: 24, 24, 24, 24
        565 => x"18151515",		-- colors: 24, 21, 21, 21
        566 => x"14141414",		-- colors: 20, 20, 20, 20
        567 => x"14151515",		-- colors: 20, 21, 21, 21
        568 => x"15161616",		-- colors: 21, 22, 22, 22
        569 => x"16151414",		-- colors: 22, 21, 20, 20
        570 => x"14141414",		-- colors: 20, 20, 20, 20
        571 => x"14141514",		-- colors: 20, 20, 21, 20
        572 => x"14141414",		-- colors: 20, 20, 20, 20
        573 => x"14141414",		-- colors: 20, 20, 20, 20
        574 => x"14141414",		-- colors: 20, 20, 20, 20

--blue car sprite


                --  sprite 0
        575 => x"27272727",		-- colors: 39, 39, 39, 39
        576 => x"27272727",		-- colors: 39, 39, 39, 39
        577 => x"27272727",		-- colors: 39, 39, 39, 39
        578 => x"27272727",		-- colors: 39, 39, 39, 39
        579 => x"27272727",		-- colors: 39, 39, 39, 39
        580 => x"27272829",		-- colors: 39, 39, 40, 41
        581 => x"28272727",		-- colors: 40, 39, 39, 39
        582 => x"27272727",		-- colors: 39, 39, 39, 39
        583 => x"27272727",		-- colors: 39, 39, 39, 39
        584 => x"2727282A",		-- colors: 39, 39, 40, 42
        585 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
        586 => x"2A2A2727",		-- colors: 42, 42, 39, 39
        587 => x"27272728",		-- colors: 39, 39, 39, 40
        588 => x"27272A2A",		-- colors: 39, 39, 42, 42
        589 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
        590 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
        591 => x"2727292D",		-- colors: 39, 39, 41, 45
        592 => x"2A2A2E2E",		-- colors: 42, 42, 46, 46
        593 => x"2E2E2E2E",		-- colors: 46, 46, 46, 46
        594 => x"2F2F2A2A",		-- colors: 47, 47, 42, 42
        595 => x"27272A2A",		-- colors: 39, 39, 42, 42
        596 => x"2E2E2E2E",		-- colors: 46, 46, 46, 46
        597 => x"2E2E2F2F",		-- colors: 46, 46, 47, 47
        598 => x"2F2F2A2A",		-- colors: 47, 47, 42, 42
        599 => x"30302E2E",		-- colors: 48, 48, 46, 46
        600 => x"2E2E2E2E",		-- colors: 46, 46, 46, 46
        601 => x"2F2F2F2F",		-- colors: 47, 47, 47, 47
        602 => x"2F2F2A2A",		-- colors: 47, 47, 42, 42
        603 => x"2A2A2E2E",		-- colors: 42, 42, 46, 46
        604 => x"2E2E2E2F",		-- colors: 46, 46, 46, 47
        605 => x"2F2F2F2F",		-- colors: 47, 47, 47, 47
        606 => x"2F2F2A2A",		-- colors: 47, 47, 42, 42
        607 => x"2A2A2E2E",		-- colors: 42, 42, 46, 46
        608 => x"2E2E2E2F",		-- colors: 46, 46, 46, 47
        609 => x"2F2F2F2F",		-- colors: 47, 47, 47, 47
        610 => x"2F2F2A2A",		-- colors: 47, 47, 42, 42
        611 => x"2A2A2E2E",		-- colors: 42, 42, 46, 46
        612 => x"2E2E2E2F",		-- colors: 46, 46, 46, 47
        613 => x"2F2F2F2F",		-- colors: 47, 47, 47, 47
        614 => x"2F2F2A2A",		-- colors: 47, 47, 42, 42
        615 => x"30302E2E",		-- colors: 48, 48, 46, 46
        616 => x"2E2E2E2E",		-- colors: 46, 46, 46, 46
        617 => x"2F2F2F2F",		-- colors: 47, 47, 47, 47
        618 => x"2F2F2A2A",		-- colors: 47, 47, 42, 42
        619 => x"27272A2A",		-- colors: 39, 39, 42, 42
        620 => x"2E2E2E2E",		-- colors: 46, 46, 46, 46
        621 => x"2E2E2F2F",		-- colors: 46, 46, 47, 47
        622 => x"2F2F2A2A",		-- colors: 47, 47, 42, 42
        623 => x"27282827",		-- colors: 39, 40, 40, 39
        624 => x"2A2A2E2E",		-- colors: 42, 42, 46, 46
        625 => x"2E2E2E2E",		-- colors: 46, 46, 46, 46
        626 => x"2F2F2A2A",		-- colors: 47, 47, 42, 42
        627 => x"27272728",		-- colors: 39, 39, 39, 40
        628 => x"29322A2A",		-- colors: 41, 50, 42, 42
        629 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
        630 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
        631 => x"27272727",		-- colors: 39, 39, 39, 39
        632 => x"2727272A",		-- colors: 39, 39, 39, 42
        633 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
        634 => x"2A2A2727",		-- colors: 42, 42, 39, 39
        635 => x"27272727",		-- colors: 39, 39, 39, 39
        636 => x"27272727",		-- colors: 39, 39, 39, 39
        637 => x"27272727",		-- colors: 39, 39, 39, 39
        638 => x"27272727",		-- colors: 39, 39, 39, 39

                --  sprite 1
        639 => x"27272727",		-- colors: 39, 39, 39, 39
        640 => x"27272727",		-- colors: 39, 39, 39, 39
        641 => x"27272727",		-- colors: 39, 39, 39, 39
        642 => x"27272727",		-- colors: 39, 39, 39, 39
        643 => x"27272727",		-- colors: 39, 39, 39, 39
        644 => x"27272929",		-- colors: 39, 39, 41, 41
        645 => x"28272727",		-- colors: 40, 39, 39, 39
        646 => x"27272727",		-- colors: 39, 39, 39, 39
        647 => x"27272728",		-- colors: 39, 39, 39, 40
        648 => x"27272A2A",		-- colors: 39, 39, 42, 42
        649 => x"2A282827",		-- colors: 42, 40, 40, 39
        650 => x"27272727",		-- colors: 39, 39, 39, 39
        651 => x"2B2B2C27",		-- colors: 43, 43, 44, 39
        652 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
        653 => x"2A2A2728",		-- colors: 42, 42, 39, 40
        654 => x"29282727",		-- colors: 41, 40, 39, 39
        655 => x"2E2E2A2A",		-- colors: 46, 46, 42, 42
        656 => x"2E2E2E2E",		-- colors: 46, 46, 46, 46
        657 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
        658 => x"2A2A2827",		-- colors: 42, 42, 40, 39
        659 => x"2E2E2A2A",		-- colors: 46, 46, 42, 42
        660 => x"2E2E2E2E",		-- colors: 46, 46, 46, 46
        661 => x"2A2A2E2E",		-- colors: 42, 42, 46, 46
        662 => x"2E2A2A28",		-- colors: 46, 42, 42, 40
        663 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
        664 => x"2A31312A",		-- colors: 42, 49, 49, 42
        665 => x"2A2A2E2E",		-- colors: 42, 42, 46, 46
        666 => x"2E2E2A2A",		-- colors: 46, 46, 42, 42
        667 => x"2E2E2E2E",		-- colors: 46, 46, 46, 46
        668 => x"2E2E2E2E",		-- colors: 46, 46, 46, 46
        669 => x"2A2A2E2E",		-- colors: 42, 42, 46, 46
        670 => x"2E2E2A2A",		-- colors: 46, 46, 42, 42
        671 => x"2A2E2E2E",		-- colors: 42, 46, 46, 46
        672 => x"2E2E2E2E",		-- colors: 46, 46, 46, 46
        673 => x"2A2A2E2E",		-- colors: 42, 42, 46, 46
        674 => x"2E2E2A2A",		-- colors: 46, 46, 42, 42
        675 => x"2E2E2E2E",		-- colors: 46, 46, 46, 46
        676 => x"2E2E2E2E",		-- colors: 46, 46, 46, 46
        677 => x"2A2A2E2E",		-- colors: 42, 42, 46, 46
        678 => x"2E2E2A2A",		-- colors: 46, 46, 42, 42
        679 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
        680 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
        681 => x"2A2A2E2E",		-- colors: 42, 42, 46, 46
        682 => x"2E2E2A2A",		-- colors: 46, 46, 42, 42
        683 => x"2E2E2A2A",		-- colors: 46, 46, 42, 42
        684 => x"2E2E2E2E",		-- colors: 46, 46, 46, 46
        685 => x"2A2A2E2E",		-- colors: 42, 42, 46, 46
        686 => x"2E2A2A28",		-- colors: 46, 42, 42, 40
        687 => x"2E2E2A2A",		-- colors: 46, 46, 42, 42
        688 => x"2E2E2E2E",		-- colors: 46, 46, 46, 46
        689 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
        690 => x"2A2A2727",		-- colors: 42, 42, 39, 39
        691 => x"33342C27",		-- colors: 51, 52, 44, 39
        692 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
        693 => x"2A2A2727",		-- colors: 42, 42, 39, 39
        694 => x"28272727",		-- colors: 40, 39, 39, 39
        695 => x"27272728",		-- colors: 39, 39, 39, 40
        696 => x"28272A2A",		-- colors: 40, 39, 42, 42
        697 => x"2A273527",		-- colors: 42, 39, 53, 39
        698 => x"27272727",		-- colors: 39, 39, 39, 39
        699 => x"27272727",		-- colors: 39, 39, 39, 39
        700 => x"27282929",		-- colors: 39, 40, 41, 41
        701 => x"29282727",		-- colors: 41, 40, 39, 39
        702 => x"27272727",		-- colors: 39, 39, 39, 39
      






       

--		****  MAP  ****
     
       
                --  sprite 0
        
                --  sprite 0
        6992 => x"07070707",		-- colors: 7, 7, 7, 7
        6993 => x"07070707",		-- colors: 7, 7, 7, 7
        6994 => x"07070707",		-- colors: 7, 7, 7, 7
        6995 => x"07070707",		-- colors: 7, 7, 7, 7
        6996 => x"07070707",		-- colors: 7, 7, 7, 7
        6997 => x"07070707",		-- colors: 7, 7, 7, 7
        6998 => x"07070707",		-- colors: 7, 7, 7, 7
        6999 => x"07070707",		-- colors: 7, 7, 7, 7
        7000 => x"07070707",		-- colors: 7, 7, 7, 7
        7001 => x"07070707",		-- colors: 7, 7, 7, 7
        7002 => x"07070707",		-- colors: 7, 7, 7, 7
        7003 => x"07070707",		-- colors: 7, 7, 7, 7
        7004 => x"07070707",		-- colors: 7, 7, 7, 7
        7005 => x"07070707",		-- colors: 7, 7, 7, 7
        7006 => x"07070707",		-- colors: 7, 7, 7, 7
        7007 => x"07070707",		-- colors: 7, 7, 7, 7
        7008 => x"07070707",		-- colors: 7, 7, 7, 7
        7009 => x"07070707",		-- colors: 7, 7, 7, 7
        7010 => x"07070707",		-- colors: 7, 7, 7, 7
        7011 => x"07070707",		-- colors: 7, 7, 7, 7
        7012 => x"07070707",		-- colors: 7, 7, 7, 7
        7013 => x"07070707",		-- colors: 7, 7, 7, 7
        7014 => x"07070707",		-- colors: 7, 7, 7, 7
        7015 => x"07070707",		-- colors: 7, 7, 7, 7
        7016 => x"07070707",		-- colors: 7, 7, 7, 7
        7017 => x"07070707",		-- colors: 7, 7, 7, 7
        7018 => x"07070707",		-- colors: 7, 7, 7, 7
        7019 => x"07070707",		-- colors: 7, 7, 7, 7
        7020 => x"07070707",		-- colors: 7, 7, 7, 7
        7021 => x"07070707",		-- colors: 7, 7, 7, 7
        7022 => x"07070707",		-- colors: 7, 7, 7, 7
        7023 => x"07070707",		-- colors: 7, 7, 7, 7
        7024 => x"07070707",		-- colors: 7, 7, 7, 7
        7025 => x"07070707",		-- colors: 7, 7, 7, 7
        7026 => x"07070707",		-- colors: 7, 7, 7, 7
        7027 => x"07070707",		-- colors: 7, 7, 7, 7
        7028 => x"07070707",		-- colors: 7, 7, 7, 7
        7029 => x"07070707",		-- colors: 7, 7, 7, 7
        7030 => x"07070707",		-- colors: 7, 7, 7, 7
        7031 => x"07070707",		-- colors: 7, 7, 7, 7
        7032 => x"07070707",		-- colors: 7, 7, 7, 7
        7033 => x"07070707",		-- colors: 7, 7, 7, 7
        7034 => x"07070707",		-- colors: 7, 7, 7, 7
        7035 => x"07070707",		-- colors: 7, 7, 7, 7
        7036 => x"07070707",		-- colors: 7, 7, 7, 7
        7037 => x"07070707",		-- colors: 7, 7, 7, 7
        7038 => x"07070707",		-- colors: 7, 7, 7, 7
        7039 => x"07070707",		-- colors: 7, 7, 7, 7
        7040 => x"07070707",		-- colors: 7, 7, 7, 7
        7041 => x"07070707",		-- colors: 7, 7, 7, 7
        7042 => x"07070707",		-- colors: 7, 7, 7, 7
        7043 => x"07070707",		-- colors: 7, 7, 7, 7
        7044 => x"07070707",		-- colors: 7, 7, 7, 7
        7045 => x"07070707",		-- colors: 7, 7, 7, 7
        7046 => x"07070707",		-- colors: 7, 7, 7, 7
        7047 => x"07070707",		-- colors: 7, 7, 7, 7
        7048 => x"07070707",		-- colors: 7, 7, 7, 7
        7049 => x"07070707",		-- colors: 7, 7, 7, 7
        7050 => x"07070707",		-- colors: 7, 7, 7, 7
        7051 => x"07070707",		-- colors: 7, 7, 7, 7
        7052 => x"07070707",		-- colors: 7, 7, 7, 7
        7053 => x"07070707",		-- colors: 7, 7, 7, 7
        7054 => x"07070707",		-- colors: 7, 7, 7, 7
        7055 => x"07070707",		-- colors: 7, 7, 7, 7

                --  sprite 1
        7056 => x"08080808",		-- colors: 8, 8, 8, 8
        7057 => x"08080808",		-- colors: 8, 8, 8, 8
        7058 => x"08080808",		-- colors: 8, 8, 8, 8
        7059 => x"08080808",		-- colors: 8, 8, 8, 8
        7060 => x"08080808",		-- colors: 8, 8, 8, 8
        7061 => x"08080808",		-- colors: 8, 8, 8, 8
        7062 => x"08080808",		-- colors: 8, 8, 8, 8
        7063 => x"08080808",		-- colors: 8, 8, 8, 8
        7064 => x"08080808",		-- colors: 8, 8, 8, 8
        7065 => x"08080808",		-- colors: 8, 8, 8, 8
        7066 => x"08080808",		-- colors: 8, 8, 8, 8
        7067 => x"08080808",		-- colors: 8, 8, 8, 8
        7068 => x"08080808",		-- colors: 8, 8, 8, 8
        7069 => x"08080808",		-- colors: 8, 8, 8, 8
        7070 => x"08080808",		-- colors: 8, 8, 8, 8
        7071 => x"08080808",		-- colors: 8, 8, 8, 8
        7072 => x"08080808",		-- colors: 8, 8, 8, 8
        7073 => x"08080808",		-- colors: 8, 8, 8, 8
        7074 => x"08080808",		-- colors: 8, 8, 8, 8
        7075 => x"08080808",		-- colors: 8, 8, 8, 8
        7076 => x"08080808",		-- colors: 8, 8, 8, 8
        7077 => x"08080808",		-- colors: 8, 8, 8, 8
        7078 => x"08080808",		-- colors: 8, 8, 8, 8
        7079 => x"08080808",		-- colors: 8, 8, 8, 8
        7080 => x"08080808",		-- colors: 8, 8, 8, 8
        7081 => x"08080808",		-- colors: 8, 8, 8, 8
        7082 => x"08080808",		-- colors: 8, 8, 8, 8
        7083 => x"08080808",		-- colors: 8, 8, 8, 8
        7084 => x"08080808",		-- colors: 8, 8, 8, 8
        7085 => x"08080808",		-- colors: 8, 8, 8, 8
        7086 => x"08080808",		-- colors: 8, 8, 8, 8
        7087 => x"08080808",		-- colors: 8, 8, 8, 8
        7088 => x"08080808",		-- colors: 8, 8, 8, 8
        7089 => x"08080808",		-- colors: 8, 8, 8, 8
        7090 => x"08080808",		-- colors: 8, 8, 8, 8
        7091 => x"08080808",		-- colors: 8, 8, 8, 8
        7092 => x"08080808",		-- colors: 8, 8, 8, 8
        7093 => x"08080808",		-- colors: 8, 8, 8, 8
        7094 => x"08080808",		-- colors: 8, 8, 8, 8
        7095 => x"08080808",		-- colors: 8, 8, 8, 8
        7096 => x"08080808",		-- colors: 8, 8, 8, 8
        7097 => x"08080808",		-- colors: 8, 8, 8, 8
        7098 => x"08080808",		-- colors: 8, 8, 8, 8
        7099 => x"08080808",		-- colors: 8, 8, 8, 8
        7100 => x"08080808",		-- colors: 8, 8, 8, 8
        7101 => x"08080808",		-- colors: 8, 8, 8, 8
        7102 => x"08080808",		-- colors: 8, 8, 8, 8
        7103 => x"08080808",		-- colors: 8, 8, 8, 8
        7104 => x"08080808",		-- colors: 8, 8, 8, 8
        7105 => x"08080808",		-- colors: 8, 8, 8, 8
        7106 => x"08080808",		-- colors: 8, 8, 8, 8
        7107 => x"08080808",		-- colors: 8, 8, 8, 8
        7108 => x"08080808",		-- colors: 8, 8, 8, 8
        7109 => x"08080808",		-- colors: 8, 8, 8, 8
        7110 => x"08080808",		-- colors: 8, 8, 8, 8
        7111 => x"08080808",		-- colors: 8, 8, 8, 8
        7112 => x"08080808",		-- colors: 8, 8, 8, 8
        7113 => x"08080808",		-- colors: 8, 8, 8, 8
        7114 => x"08080808",		-- colors: 8, 8, 8, 8
        7115 => x"08080808",		-- colors: 8, 8, 8, 8
        7116 => x"08080808",		-- colors: 8, 8, 8, 8
        7117 => x"08080808",		-- colors: 8, 8, 8, 8
        7118 => x"08080808",		-- colors: 8, 8, 8, 8
        7119 => x"08080808",		-- colors: 8, 8, 8, 8

                --  sprite 2
        7120 => x"09090909",		-- colors: 9, 9, 9, 9
        7121 => x"09090909",		-- colors: 9, 9, 9, 9
        7122 => x"09090909",		-- colors: 9, 9, 9, 9
        7123 => x"09090909",		-- colors: 9, 9, 9, 9
        7124 => x"09090909",		-- colors: 9, 9, 9, 9
        7125 => x"09090909",		-- colors: 9, 9, 9, 9
        7126 => x"09090909",		-- colors: 9, 9, 9, 9
        7127 => x"09090909",		-- colors: 9, 9, 9, 9
        7128 => x"09090909",		-- colors: 9, 9, 9, 9
        7129 => x"09090909",		-- colors: 9, 9, 9, 9
        7130 => x"09090909",		-- colors: 9, 9, 9, 9
        7131 => x"09090909",		-- colors: 9, 9, 9, 9
        7132 => x"09090909",		-- colors: 9, 9, 9, 9
        7133 => x"09090909",		-- colors: 9, 9, 9, 9
        7134 => x"09090909",		-- colors: 9, 9, 9, 9
        7135 => x"09090909",		-- colors: 9, 9, 9, 9
        7136 => x"09090909",		-- colors: 9, 9, 9, 9
        7137 => x"09090909",		-- colors: 9, 9, 9, 9
        7138 => x"09090909",		-- colors: 9, 9, 9, 9
        7139 => x"09090909",		-- colors: 9, 9, 9, 9
        7140 => x"09090909",		-- colors: 9, 9, 9, 9
        7141 => x"09090909",		-- colors: 9, 9, 9, 9
        7142 => x"09090909",		-- colors: 9, 9, 9, 9
        7143 => x"09090909",		-- colors: 9, 9, 9, 9
        7144 => x"09090909",		-- colors: 9, 9, 9, 9
        7145 => x"09090909",		-- colors: 9, 9, 9, 9
        7146 => x"09090909",		-- colors: 9, 9, 9, 9
        7147 => x"09090909",		-- colors: 9, 9, 9, 9
        7148 => x"09090909",		-- colors: 9, 9, 9, 9
        7149 => x"09090909",		-- colors: 9, 9, 9, 9
        7150 => x"09090909",		-- colors: 9, 9, 9, 9
        7151 => x"09090909",		-- colors: 9, 9, 9, 9
        7152 => x"09090909",		-- colors: 9, 9, 9, 9
        7153 => x"09090909",		-- colors: 9, 9, 9, 9
        7154 => x"09090909",		-- colors: 9, 9, 9, 9
        7155 => x"09090909",		-- colors: 9, 9, 9, 9
        7156 => x"09090909",		-- colors: 9, 9, 9, 9
        7157 => x"09090909",		-- colors: 9, 9, 9, 9
        7158 => x"09090909",		-- colors: 9, 9, 9, 9
        7159 => x"09090909",		-- colors: 9, 9, 9, 9
        7160 => x"09090909",		-- colors: 9, 9, 9, 9
        7161 => x"09090909",		-- colors: 9, 9, 9, 9
        7162 => x"09090909",		-- colors: 9, 9, 9, 9
        7163 => x"09090909",		-- colors: 9, 9, 9, 9
        7164 => x"09090909",		-- colors: 9, 9, 9, 9
        7165 => x"09090909",		-- colors: 9, 9, 9, 9
        7166 => x"09090909",		-- colors: 9, 9, 9, 9
        7167 => x"09090909",		-- colors: 9, 9, 9, 9
        7168 => x"09090909",		-- colors: 9, 9, 9, 9
        7169 => x"09090909",		-- colors: 9, 9, 9, 9
        7170 => x"09090909",		-- colors: 9, 9, 9, 9
        7171 => x"09090909",		-- colors: 9, 9, 9, 9
        7172 => x"09090909",		-- colors: 9, 9, 9, 9
        7173 => x"09090909",		-- colors: 9, 9, 9, 9
        7174 => x"09090909",		-- colors: 9, 9, 9, 9
        7175 => x"09090909",		-- colors: 9, 9, 9, 9
        7176 => x"09090909",		-- colors: 9, 9, 9, 9
        7177 => x"09090909",		-- colors: 9, 9, 9, 9
        7178 => x"09090909",		-- colors: 9, 9, 9, 9
        7179 => x"09090909",		-- colors: 9, 9, 9, 9
        7180 => x"09090909",		-- colors: 9, 9, 9, 9
        7181 => x"09090909",		-- colors: 9, 9, 9, 9
        7182 => x"09090909",		-- colors: 9, 9, 9, 9
        7183 => x"09090909",		-- colors: 9, 9, 9, 9

                --  sprite 3
        7184 => x"0A0A0A0A",		-- colors: 10, 10, 10, 10
        7185 => x"0A0A0A0A",		-- colors: 10, 10, 10, 10
        7186 => x"0A0A0A0A",		-- colors: 10, 10, 10, 10
        7187 => x"0A0A0A0A",		-- colors: 10, 10, 10, 10
        7188 => x"0A0A0A0A",		-- colors: 10, 10, 10, 10
        7189 => x"0A0A0A0A",		-- colors: 10, 10, 10, 10
        7190 => x"0A0A0A0A",		-- colors: 10, 10, 10, 10
        7191 => x"0A0A0A0A",		-- colors: 10, 10, 10, 10
        7192 => x"0A0A0A0A",		-- colors: 10, 10, 10, 10
        7193 => x"0A0A0A0A",		-- colors: 10, 10, 10, 10
        7194 => x"0A0A0A0A",		-- colors: 10, 10, 10, 10
        7195 => x"0A0A0A0A",		-- colors: 10, 10, 10, 10
        7196 => x"0A0A0A0A",		-- colors: 10, 10, 10, 10
        7197 => x"0A0A0A0A",		-- colors: 10, 10, 10, 10
        7198 => x"0A0A0A0A",		-- colors: 10, 10, 10, 10
        7199 => x"0A0A0A0A",		-- colors: 10, 10, 10, 10
        7200 => x"0A0A0A0A",		-- colors: 10, 10, 10, 10
        7201 => x"0A0A0A0A",		-- colors: 10, 10, 10, 10
        7202 => x"0A0A0A0A",		-- colors: 10, 10, 10, 10
        7203 => x"0A0A0A0A",		-- colors: 10, 10, 10, 10
        7204 => x"0A0A0A0A",		-- colors: 10, 10, 10, 10
        7205 => x"0A0A0A0A",		-- colors: 10, 10, 10, 10
        7206 => x"0A0A0A0A",		-- colors: 10, 10, 10, 10
        7207 => x"0A0A0A0A",		-- colors: 10, 10, 10, 10
        7208 => x"0A0A0A0A",		-- colors: 10, 10, 10, 10
        7209 => x"0A0A0A0A",		-- colors: 10, 10, 10, 10
        7210 => x"0A0A0A0A",		-- colors: 10, 10, 10, 10
        7211 => x"0A0A0A0A",		-- colors: 10, 10, 10, 10
        7212 => x"0A0A0A0A",		-- colors: 10, 10, 10, 10
        7213 => x"0A0A0A0A",		-- colors: 10, 10, 10, 10
        7214 => x"0A0A0A0A",		-- colors: 10, 10, 10, 10
        7215 => x"0A0A0A0A",		-- colors: 10, 10, 10, 10
        7216 => x"0A0A0A0A",		-- colors: 10, 10, 10, 10
        7217 => x"0A0A0A0A",		-- colors: 10, 10, 10, 10
        7218 => x"0A0A0A0A",		-- colors: 10, 10, 10, 10
        7219 => x"0A0A0A0A",		-- colors: 10, 10, 10, 10
        7220 => x"0A0A0A0A",		-- colors: 10, 10, 10, 10
        7221 => x"0A0A0A0A",		-- colors: 10, 10, 10, 10
        7222 => x"0A0A0A0A",		-- colors: 10, 10, 10, 10
        7223 => x"0A0A0A0A",		-- colors: 10, 10, 10, 10
        7224 => x"0A0A0A0A",		-- colors: 10, 10, 10, 10
        7225 => x"0A0A0A0A",		-- colors: 10, 10, 10, 10
        7226 => x"0A0A0A0A",		-- colors: 10, 10, 10, 10
        7227 => x"0A0A0A0A",		-- colors: 10, 10, 10, 10
        7228 => x"0A0A0A0A",		-- colors: 10, 10, 10, 10
        7229 => x"0A0A0A0A",		-- colors: 10, 10, 10, 10
        7230 => x"0A0A0A0A",		-- colors: 10, 10, 10, 10
        7231 => x"0A0A0A0A",		-- colors: 10, 10, 10, 10
        7232 => x"0A0A0A0A",		-- colors: 10, 10, 10, 10
        7233 => x"0A0A0A0A",		-- colors: 10, 10, 10, 10
        7234 => x"0A0A0A0A",		-- colors: 10, 10, 10, 10
        7235 => x"0A0A0A0A",		-- colors: 10, 10, 10, 10
        7236 => x"0A0A0A0A",		-- colors: 10, 10, 10, 10
        7237 => x"0A0A0A0A",		-- colors: 10, 10, 10, 10
        7238 => x"0A0A0A0A",		-- colors: 10, 10, 10, 10
        7239 => x"0A0A0A0A",		-- colors: 10, 10, 10, 10
        7240 => x"0A0A0A0A",		-- colors: 10, 10, 10, 10
        7241 => x"0A0A0A0A",		-- colors: 10, 10, 10, 10
        7242 => x"0A0A0A0A",		-- colors: 10, 10, 10, 10
        7243 => x"0A0A0A0A",		-- colors: 10, 10, 10, 10
        7244 => x"0A0A0A0A",		-- colors: 10, 10, 10, 10
        7245 => x"0A0A0A0A",		-- colors: 10, 10, 10, 10
        7246 => x"0A0A0A0A",		-- colors: 10, 10, 10, 10
        7247 => x"0A0A0A0A",		-- colors: 10, 10, 10, 10

                --  sprite 4
        7248 => x"0B0B0B0B",		-- colors: 11, 11, 11, 11
        7249 => x"0B0B0C0B",		-- colors: 11, 11, 12, 11
        7250 => x"0C0D0B0B",		-- colors: 12, 13, 11, 11
        7251 => x"0B0B0B0B",		-- colors: 11, 11, 11, 11
        7252 => x"0B0B0B0C",		-- colors: 11, 11, 11, 12
        7253 => x"0C0C0C0C",		-- colors: 12, 12, 12, 12
        7254 => x"0C0C0C0C",		-- colors: 12, 12, 12, 12
        7255 => x"0B0B0B0B",		-- colors: 11, 11, 11, 11
        7256 => x"0B0B0C0C",		-- colors: 11, 11, 12, 12
        7257 => x"0C0C0E0C",		-- colors: 12, 12, 14, 12
        7258 => x"0C0C0C0C",		-- colors: 12, 12, 12, 12
        7259 => x"0C0B0B0B",		-- colors: 12, 11, 11, 11
        7260 => x"0B0B0C0C",		-- colors: 11, 11, 12, 12
        7261 => x"0C0C0C0C",		-- colors: 12, 12, 12, 12
        7262 => x"0C0C0C0F",		-- colors: 12, 12, 12, 15
        7263 => x"0C0C0B0B",		-- colors: 12, 12, 11, 11
        7264 => x"0B0B0B0C",		-- colors: 11, 11, 11, 12
        7265 => x"0C0C0C0C",		-- colors: 12, 12, 12, 12
        7266 => x"0C0C0C0C",		-- colors: 12, 12, 12, 12
        7267 => x"0C0C0C0B",		-- colors: 12, 12, 12, 11
        7268 => x"0B0B0C0C",		-- colors: 11, 11, 12, 12
        7269 => x"0C0C0C0C",		-- colors: 12, 12, 12, 12
        7270 => x"0C0C0C0C",		-- colors: 12, 12, 12, 12
        7271 => x"0C0C0C0B",		-- colors: 12, 12, 12, 11
        7272 => x"0B0C0C0C",		-- colors: 11, 12, 12, 12
        7273 => x"0C0C0C0C",		-- colors: 12, 12, 12, 12
        7274 => x"0C0C0C0C",		-- colors: 12, 12, 12, 12
        7275 => x"0C0C0B0B",		-- colors: 12, 12, 11, 11
        7276 => x"0B0C0C0C",		-- colors: 11, 12, 12, 12
        7277 => x"0C0C0C0C",		-- colors: 12, 12, 12, 12
        7278 => x"0C100C0C",		-- colors: 12, 16, 12, 12
        7279 => x"0C0C0B0B",		-- colors: 12, 12, 11, 11
        7280 => x"0B0C0C0C",		-- colors: 11, 12, 12, 12
        7281 => x"0C0C0E11",		-- colors: 12, 12, 14, 17
        7282 => x"110C0C0C",		-- colors: 17, 12, 12, 12
        7283 => x"0C0C0B0B",		-- colors: 12, 12, 11, 11
        7284 => x"0B0B0C0C",		-- colors: 11, 11, 12, 12
        7285 => x"0C0E0C11",		-- colors: 12, 14, 12, 17
        7286 => x"110C0C0C",		-- colors: 17, 12, 12, 12
        7287 => x"0C0C0B0B",		-- colors: 12, 12, 11, 11
        7288 => x"0B0B0C0C",		-- colors: 11, 11, 12, 12
        7289 => x"0C0C0C0C",		-- colors: 12, 12, 12, 12
        7290 => x"0C0C0C0C",		-- colors: 12, 12, 12, 12
        7291 => x"0B0B0B0B",		-- colors: 11, 11, 11, 11
        7292 => x"0B0B0C0C",		-- colors: 11, 11, 12, 12
        7293 => x"0C0C0C0C",		-- colors: 12, 12, 12, 12
        7294 => x"0C0C0C0B",		-- colors: 12, 12, 12, 11
        7295 => x"0B0B0B0B",		-- colors: 11, 11, 11, 11
        7296 => x"0B0B0C0C",		-- colors: 11, 11, 12, 12
        7297 => x"0C0C0C0C",		-- colors: 12, 12, 12, 12
        7298 => x"0C0C0C0B",		-- colors: 12, 12, 12, 11
        7299 => x"0B0B0B0B",		-- colors: 11, 11, 11, 11
        7300 => x"0B0B0B0C",		-- colors: 11, 11, 11, 12
        7301 => x"0B0B0C0C",		-- colors: 11, 11, 12, 12
        7302 => x"0C0C0B0B",		-- colors: 12, 12, 11, 11
        7303 => x"0B0B0B0B",		-- colors: 11, 11, 11, 11
        7304 => x"0B0B0B0B",		-- colors: 11, 11, 11, 11
        7305 => x"0B0B0C0C",		-- colors: 11, 11, 12, 12
        7306 => x"0C0B0B0B",		-- colors: 12, 11, 11, 11
        7307 => x"0B0B0B0B",		-- colors: 11, 11, 11, 11
        7308 => x"0B0B0B0B",		-- colors: 11, 11, 11, 11
        7309 => x"0B0B0B0B",		-- colors: 11, 11, 11, 11
        7310 => x"0B0B0B0B",		-- colors: 11, 11, 11, 11
        7311 => x"0B0B0B0B",		-- colors: 11, 11, 11, 11
others => x"00000000"
	);


begin

	process(i_clk)
	begin
		if rising_edge(i_clk) then
			-- memory write --
			if i_we = '1' then
				mem(to_integer(unsigned(i_w_addr))) <= i_data;
			end if;
			-- memory read -- 
			o_data <= mem(to_integer(unsigned(i_r_addr)));
			
		end if; 
	end process;

end architecture arch;
