
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity ram is
	generic
	(
		DATA_WIDTH : natural := 32;		    -- 4 byte one line of memory
		ADDR_WIDTH : natural := 13			    -- 24576 bytes size of memory
	);

	port(
		i_clk    : in  std_logic;
		i_r_addr : in  std_logic_vector(ADDR_WIDTH-1 downto 0);
		i_data   : in  std_logic_vector(DATA_WIDTH-1 downto 0);
		i_we     : in  std_logic;
		i_w_addr : in  std_logic_vector(ADDR_WIDTH-1 downto 0);
		o_data   : out std_logic_vector(DATA_WIDTH-1 downto 0)
	);
end entity ram;

architecture arch of ram is

	type ram_t is array (0 to 2**ADDR_WIDTH-1) of std_logic_vector(DATA_WIDTH-1 downto 0);


-- GENERATED BY BC_MEM_PACKER

-- DATE: Thu May 18 16:01:02 2017

	signal mem : ram_t := (

--			***** COLOR PALLETE *****

		-- fellas
		--0 =>	x"000C4CC8", 
		--1 =>	x"00A8D8FC", 
		--2 =>	x"00000000", 
		--3 =>	x"00EC3820", 
		--4 =>	x"0000A800", 
		--5 =>	x"00FCFCFC", 
		--6 =>	x"00747474",
		--7 =>	x"00C0C0C0",


--kirby colors
        8 0x"00000000",
        9 0x"00ea8bff",
        10 0x"00e98afe",
        11 0x"003d3d40",
        12 0x"00811699",
        13 0x"00ea8aff",
        14 0x"000303d5",
--trava colors
	35=> x"00353b39",
	36=> x"000cac83",
	37=> x"00ffffff",
	38=> x"009b6f2e",
	39=> x"00000000",
	40=> x"0019704d",
	41=> x"00010101",
	42=> x"001b714d",
	43=> x"001b714e",
	44=> x"001c714e",
	45=> x"001a6e4f",
	
--deblo
	46 0x"00000000
        47 0x"0008072c
        
--blue_car

          48 => 0x"0000000000"
          49 => 0x"0000000001"
          50 => 0x"0000000002"
          51 => 0x"000008072c"
          52 => 0x"0000070102"
          53 => 0x"0000020102"
          54 => 0x"0000010002"
          55 => 0x"0000ab1c2b"
          56 => 0x"0000b09256"
          57 => 0x"00000a072b"
          58 => 0x"000007062b"
          59 => 0x"0000aa1b2c"
          60 => 0x"000000dcd6"
          61 => 0x"000016092c"
          62 => 0x"000019092c"
          63 => 0x"000012082c"
          64 => 0x"0000a81b2e"
          65 => 0x"0000a81b32"
          66 => 0x"0000a81b2f"
          67 => 0x"0000a91c2c"
          68 => 0x"0000b09156"
          69 => 0x"0000b19357"
          70 => 0x"0000010106"
          71 => 0x"000007072c"
          72 => 0x"0000020101"
          73 => 0x"0000010000"
          74 => 0x"0000060102"
          75 => 0x"0000010102"
        
--
	
	
	

	        --  heart colors	
        --57 => 	x"00000000",
        --58 => 	x"002131b5",
        --59 =>	x"00c4cdfe",
            -- orange and red for grandpa and rupees
        --60 =>   x"003b9bff", -- orange 
	--	61 =>	x"00002bdb", -- red

	--	62 =>	x"003C9AFC", -- Unused
	--	63 =>	x"003199FF", -- Unused

            --  ADDED SPRITES HERE
          -- RUPEE SPRITE
		64 => x"0202020F",
		65 => x"3C020202",
		66 => x"02020202",
		67 => x"02020202",
		68 => x"02020F0F",
		69 => x"3C3C0202",
		70 => x"02020202",
		71 => x"02020202",
		72 => x"020F0F0F",
		73 => x"3C3C3C02",
		74 => x"02020202",
		75 => x"02020202",
		76 => x"0F3C0F3C",
		77 => x"023C023C",
		78 => x"02020202",
		79 => x"02020202",
		80 => x"0F0F3C3C",
		81 => x"3C023C3C",
		82 => x"02020202",
		83 => x"02020202",
		84 => x"0F0F3C3C",
		85 => x"3C023C3C",
		86 => x"02020202",
		87 => x"02020202",
		88 => x"0F0F3C3C",
		89 => x"3C023C3C",
		90 => x"02020202",
		91 => x"02020202",
		92 => x"0F0F3C3C",
		93 => x"3C023C3C",
		94 => x"02020202",
		95 => x"02020202",
		96 => x"0F0F3C3C",
		97 => x"3C023C3C",
		98 => x"02020202",
		99 => x"02020202",
		100 => x"0F0F3C3C",
		101 => x"3C023C3C",
		102 => x"02020202",
		103 => x"02020202",
		104 => x"0F0F3C3C",
		105 => x"3C023C3C",
		106 => x"02020202",
		107 => x"02020202",
		108 => x"0F3C0F3C",
		109 => x"3C023C3C",
		110 => x"02020202",
		111 => x"02020202",
		112 => x"3C3C3C0F",
		113 => x"023C023C",
		114 => x"02020202",
		115 => x"02020202",
		116 => x"023C3C3C",
		117 => x"3C3C3C02",
		118 => x"02020202",
		119 => x"02020202",
		120 => x"02023C3C",
		121 => x"3C3C0202",
		122 => x"02020202",
		123 => x"02020202",
		124 => x"0202023C",
		125 => x"3C020202",
		126 => x"02020202",
		127 => x"02020202",

          -- BOMB SPRITE
		128 => x"02020202",
		129 => x"020F0202",
		130 => x"02020202",
		131 => x"02020202",
		132 => x"02020202",
		133 => x"020F0202",
		134 => x"02020202",
		135 => x"02020202",
		136 => x"02020202",
		137 => x"02020F02",
		138 => x"02020202",
		139 => x"02020202",
		140 => x"02020202",
		141 => x"0202020F",
		142 => x"02020202",
		143 => x"02020202",
		144 => x"02020202",
		145 => x"0202020F",
		146 => x"02020202",
		147 => x"02020202",
		148 => x"02020202",
		149 => x"02020F02",
		150 => x"02020202",
		151 => x"02020202",
		152 => x"02020D0D",
		153 => x"0D0D0202",
		154 => x"02020202",
		155 => x"02020202",
		156 => x"020D2E2E",
		157 => x"0D0D0D02",
		158 => x"02020202",
		159 => x"02020202",
		160 => x"0D2E0F2E",
		161 => x"0D0D0D0D",
		162 => x"02020202",
		163 => x"02020202",
		164 => x"0D2E2E0D",
		165 => x"0D0D0D0D",
		166 => x"02020202",
		167 => x"02020202",
		168 => x"0D0D0D0D",
		169 => x"0D0D0D0D",
		170 => x"02020202",
		171 => x"02020202",
		172 => x"0D0D0D0D",
		173 => x"0D0D0D0D",
		174 => x"02020202",
		175 => x"02020202",
		176 => x"020D0D0D",
		177 => x"0D0D0D02",
		178 => x"02020202",
		179 => x"02020202",
		180 => x"02020D0D",
		181 => x"0D0D0202",
		182 => x"02020202",
		183 => x"02020202",
		184 => x"02020202",
		185 => x"02020202",
		186 => x"02020202",
		187 => x"02020202",
		188 => x"02020202",
		189 => x"02020202",
		190 => x"02020202",
		191 => x"02020202",

--			***** 16x16 IMAGES *****
--			OVERWORLD SPRITES
        
        --kirby sprites        
               
                --  sprite 0
        255 => x"08080808",		-- colors: 8, 8, 8, 8
        256 => x"08080808",		-- colors: 8, 8, 8, 8
        257 => x"08080808",		-- colors: 8, 8, 8, 8
        258 => x"08080808",		-- colors: 8, 8, 8, 8
        259 => x"08080808",		-- colors: 8, 8, 8, 8
        260 => x"08080808",		-- colors: 8, 8, 8, 8
        261 => x"08080808",		-- colors: 8, 8, 8, 8
        262 => x"08080808",		-- colors: 8, 8, 8, 8
        263 => x"08080808",		-- colors: 8, 8, 8, 8
        264 => x"08080808",		-- colors: 8, 8, 8, 8
        265 => x"08080808",		-- colors: 8, 8, 8, 8
        266 => x"08080808",		-- colors: 8, 8, 8, 8
        267 => x"08080808",		-- colors: 8, 8, 8, 8
        268 => x"08080808",		-- colors: 8, 8, 8, 8
        269 => x"08080808",		-- colors: 8, 8, 8, 8
        270 => x"08080808",		-- colors: 8, 8, 8, 8
        271 => x"08080808",		-- colors: 8, 8, 8, 8
        272 => x"08080808",		-- colors: 8, 8, 8, 8
        273 => x"08080808",		-- colors: 8, 8, 8, 8
        274 => x"08080808",		-- colors: 8, 8, 8, 8
        275 => x"08080808",		-- colors: 8, 8, 8, 8
        276 => x"08080808",		-- colors: 8, 8, 8, 8
        277 => x"08080808",		-- colors: 8, 8, 8, 8
        278 => x"08080808",		-- colors: 8, 8, 8, 8
        279 => x"08080808",		-- colors: 8, 8, 8, 8
        280 => x"08080808",		-- colors: 8, 8, 8, 8
        281 => x"08080808",		-- colors: 8, 8, 8, 8
        282 => x"08080808",		-- colors: 8, 8, 8, 8
        283 => x"08080808",		-- colors: 8, 8, 8, 8
        284 => x"08080909",		-- colors: 8, 8, 9, 9
        285 => x"090A0808",		-- colors: 9, 10, 8, 8
        286 => x"08080808",		-- colors: 8, 8, 8, 8
        287 => x"08080808",		-- colors: 8, 8, 8, 8
        288 => x"08090909",		-- colors: 8, 9, 9, 9
        289 => x"09090908",		-- colors: 9, 9, 9, 8
        290 => x"08080808",		-- colors: 8, 8, 8, 8
        291 => x"08080808",		-- colors: 8, 8, 8, 8
        292 => x"09090B09",		-- colors: 9, 9, 11, 9
        293 => x"090B0909",		-- colors: 9, 11, 9, 9
        294 => x"08080808",		-- colors: 8, 8, 8, 8
        295 => x"08080809",		-- colors: 8, 8, 8, 9
        296 => x"09090B09",		-- colors: 9, 9, 11, 9
        297 => x"090B0909",		-- colors: 9, 11, 9, 9
        298 => x"09080808",		-- colors: 9, 8, 8, 8
        299 => x"08080809",		-- colors: 8, 8, 8, 9
        300 => x"090C0909",		-- colors: 9, 12, 9, 9
        301 => x"09090C09",		-- colors: 9, 9, 12, 9
        302 => x"09080808",		-- colors: 9, 8, 8, 8
        303 => x"08080808",		-- colors: 8, 8, 8, 8
        304 => x"0D090909",		-- colors: 13, 9, 9, 9
        305 => x"09090909",		-- colors: 9, 9, 9, 9
        306 => x"08080808",		-- colors: 8, 8, 8, 8
        307 => x"08080808",		-- colors: 8, 8, 8, 8
        308 => x"08090909",		-- colors: 8, 9, 9, 9
        309 => x"09090908",		-- colors: 9, 9, 9, 8
        310 => x"08080808",		-- colors: 8, 8, 8, 8
        311 => x"08080808",		-- colors: 8, 8, 8, 8
        312 => x"08080909",		-- colors: 8, 8, 9, 9
        313 => x"09090808",		-- colors: 9, 9, 8, 8
        314 => x"08080808",		-- colors: 8, 8, 8, 8
        315 => x"08080808",		-- colors: 8, 8, 8, 8
        316 => x"080E0E08",		-- colors: 8, 14, 14, 8
        317 => x"080E0E08",		-- colors: 8, 14, 14, 8
        318 => x"08080808",		-- colors: 8, 8, 8, 8
        
        --deblo sprite
        
                --  sprite 0
        319 => x"2E2E2E2E",		-- colors: 46, 46, 46, 46
        320 => x"2E2E2E2E",		-- colors: 46, 46, 46, 46
        321 => x"2E2E2E2E",		-- colors: 46, 46, 46, 46
        322 => x"2E2E2E2E",		-- colors: 46, 46, 46, 46
        323 => x"2E2E2E2E",		-- colors: 46, 46, 46, 46
        324 => x"2E2E2E2E",		-- colors: 46, 46, 46, 46
        325 => x"2E2E2E2E",		-- colors: 46, 46, 46, 46
        326 => x"2E2E2E2E",		-- colors: 46, 46, 46, 46
        327 => x"2E2E2E2E",		-- colors: 46, 46, 46, 46
        328 => x"2E2E2E2E",		-- colors: 46, 46, 46, 46
        329 => x"2E2E2E2E",		-- colors: 46, 46, 46, 46
        330 => x"2E2E2E2E",		-- colors: 46, 46, 46, 46
        331 => x"2E2E2E2E",		-- colors: 46, 46, 46, 46
        332 => x"2E2E2E2E",		-- colors: 46, 46, 46, 46
        333 => x"2E2E2E2E",		-- colors: 46, 46, 46, 46
        334 => x"2E2E2E2E",		-- colors: 46, 46, 46, 46
        335 => x"2E2E2E2E",		-- colors: 46, 46, 46, 46
        336 => x"2E2E2E2E",		-- colors: 46, 46, 46, 46
        337 => x"2E2E2E2E",		-- colors: 46, 46, 46, 46
        338 => x"2E2E2E2E",		-- colors: 46, 46, 46, 46
        339 => x"2E2E2E2E",		-- colors: 46, 46, 46, 46
        340 => x"2E2E2E2E",		-- colors: 46, 46, 46, 46
        341 => x"2E2E2E2E",		-- colors: 46, 46, 46, 46
        342 => x"2E2E2E2E",		-- colors: 46, 46, 46, 46
        343 => x"2E2E2E2E",		-- colors: 46, 46, 46, 46
        344 => x"2E2E2E2E",		-- colors: 46, 46, 46, 46
        345 => x"2E2E2E2E",		-- colors: 46, 46, 46, 46
        346 => x"2E2E2E2E",		-- colors: 46, 46, 46, 46
        347 => x"2F2F2F2F",		-- colors: 47, 47, 47, 47
        348 => x"2F2F2F2F",		-- colors: 47, 47, 47, 47
        349 => x"2F2F2F2F",		-- colors: 47, 47, 47, 47
        350 => x"2F2F2F2F",		-- colors: 47, 47, 47, 47
        351 => x"2F2F2F2F",		-- colors: 47, 47, 47, 47
        352 => x"2F2F2F2F",		-- colors: 47, 47, 47, 47
        353 => x"2F2F2F2F",		-- colors: 47, 47, 47, 47
        354 => x"2F2F2F2F",		-- colors: 47, 47, 47, 47
        355 => x"2F2F2F2F",		-- colors: 47, 47, 47, 47
        356 => x"2F2F2F2F",		-- colors: 47, 47, 47, 47
        357 => x"2F2F2F2F",		-- colors: 47, 47, 47, 47
        358 => x"2F2F2F2F",		-- colors: 47, 47, 47, 47
        359 => x"2F2F2F2F",		-- colors: 47, 47, 47, 47
        360 => x"2F2F2F2F",		-- colors: 47, 47, 47, 47
        361 => x"2F2F2F2F",		-- colors: 47, 47, 47, 47
        362 => x"2F2F2F2F",		-- colors: 47, 47, 47, 47
        363 => x"2F2F2F2F",		-- colors: 47, 47, 47, 47
        364 => x"2F2F2F2F",		-- colors: 47, 47, 47, 47
        365 => x"2F2F2F2F",		-- colors: 47, 47, 47, 47
        366 => x"2F2F2F2F",		-- colors: 47, 47, 47, 47
        367 => x"2F2F2F2F",		-- colors: 47, 47, 47, 47
        368 => x"2F2F2F2F",		-- colors: 47, 47, 47, 47
        369 => x"2F2F2F2F",		-- colors: 47, 47, 47, 47
        370 => x"2F2F2F2F",		-- colors: 47, 47, 47, 47
        371 => x"2F2F2F2F",		-- colors: 47, 47, 47, 47
        372 => x"2F2F2F2F",		-- colors: 47, 47, 47, 47
        373 => x"2F2F2F2F",		-- colors: 47, 47, 47, 47
        374 => x"2F2F2F2F",		-- colors: 47, 47, 47, 47
        375 => x"2F2F2F2F",		-- colors: 47, 47, 47, 47
        376 => x"2F2F2F2F",		-- colors: 47, 47, 47, 47
        377 => x"2F2F2F2F",		-- colors: 47, 47, 47, 47
        378 => x"2F2F2F2F",		-- colors: 47, 47, 47, 47
        379 => x"2F2F2F2F",		-- colors: 47, 47, 47, 47
        380 => x"2F2F2F2F",		-- colors: 47, 47, 47, 47
        381 => x"2F2F2F2F",		-- colors: 47, 47, 47, 47
        382 => x"2F2F2F2F",		-- colors: 47, 47, 47, 47

                --  sprite 1
        383 => x"2E2E2E2E",		-- colors: 46, 46, 46, 46
        384 => x"2E2E2E2E",		-- colors: 46, 46, 46, 46
        385 => x"2E2E2E2E",		-- colors: 46, 46, 46, 46
        386 => x"2E2E2E2E",		-- colors: 46, 46, 46, 46
        387 => x"2E2E2E2E",		-- colors: 46, 46, 46, 46
        388 => x"2E2E2E2E",		-- colors: 46, 46, 46, 46
        389 => x"2E2E2E2E",		-- colors: 46, 46, 46, 46
        390 => x"2E2E2E2E",		-- colors: 46, 46, 46, 46
        391 => x"2E2E2E2E",		-- colors: 46, 46, 46, 46
        392 => x"2E2E2E2E",		-- colors: 46, 46, 46, 46
        393 => x"2E2E2E2E",		-- colors: 46, 46, 46, 46
        394 => x"2E2E2E2E",		-- colors: 46, 46, 46, 46
        395 => x"2E2E2E2E",		-- colors: 46, 46, 46, 46
        396 => x"2E2E2E2E",		-- colors: 46, 46, 46, 46
        397 => x"2E2E2E2E",		-- colors: 46, 46, 46, 46
        398 => x"2E2E2E2E",		-- colors: 46, 46, 46, 46
        399 => x"2E2E2E2E",		-- colors: 46, 46, 46, 46
        400 => x"2E2E2E2E",		-- colors: 46, 46, 46, 46
        401 => x"2E2E2E2E",		-- colors: 46, 46, 46, 46
        402 => x"2E2E2E2E",		-- colors: 46, 46, 46, 46
        403 => x"2E2E2E2E",		-- colors: 46, 46, 46, 46
        404 => x"2E2E2E2E",		-- colors: 46, 46, 46, 46
        405 => x"2E2E2E2E",		-- colors: 46, 46, 46, 46
        406 => x"2E2E2E2E",		-- colors: 46, 46, 46, 46
        407 => x"2E2E2E2E",		-- colors: 46, 46, 46, 46
        408 => x"2E2E2E2E",		-- colors: 46, 46, 46, 46
        409 => x"2E2E2E2E",		-- colors: 46, 46, 46, 46
        410 => x"2E2E2E2E",		-- colors: 46, 46, 46, 46
        411 => x"2F2F2F2F",		-- colors: 47, 47, 47, 47
        412 => x"2F2F2F2F",		-- colors: 47, 47, 47, 47
        413 => x"2F2F2F2F",		-- colors: 47, 47, 47, 47
        414 => x"2F2F2F2F",		-- colors: 47, 47, 47, 47
        415 => x"2F2F2F2F",		-- colors: 47, 47, 47, 47
        416 => x"2F2F2F2F",		-- colors: 47, 47, 47, 47
        417 => x"2F2F2F2F",		-- colors: 47, 47, 47, 47
        418 => x"2F2F2F2F",		-- colors: 47, 47, 47, 47
        419 => x"2F2F2F2F",		-- colors: 47, 47, 47, 47
        420 => x"2F2F2F2F",		-- colors: 47, 47, 47, 47
        421 => x"2F2F2F2F",		-- colors: 47, 47, 47, 47
        422 => x"2F2F2F2F",		-- colors: 47, 47, 47, 47
        423 => x"2F2F2F2F",		-- colors: 47, 47, 47, 47
        424 => x"2F2F2F2F",		-- colors: 47, 47, 47, 47
        425 => x"2F2F2F2F",		-- colors: 47, 47, 47, 47
        426 => x"2F2F2F2F",		-- colors: 47, 47, 47, 47
        427 => x"2F2F2F2F",		-- colors: 47, 47, 47, 47
        428 => x"2F2F2F2F",		-- colors: 47, 47, 47, 47
        429 => x"2F2F2F2F",		-- colors: 47, 47, 47, 47
        430 => x"2F2F2F2F",		-- colors: 47, 47, 47, 47
        431 => x"2F2F2F2F",		-- colors: 47, 47, 47, 47
        432 => x"2F2F2F2F",		-- colors: 47, 47, 47, 47
        433 => x"2F2F2F2F",		-- colors: 47, 47, 47, 47
        434 => x"2F2F2F2F",		-- colors: 47, 47, 47, 47
        435 => x"2F2F2F2F",		-- colors: 47, 47, 47, 47
        436 => x"2F2F2F2F",		-- colors: 47, 47, 47, 47
        437 => x"2F2F2F2F",		-- colors: 47, 47, 47, 47
        438 => x"2F2F2F2F",		-- colors: 47, 47, 47, 47
        439 => x"2F2F2F2F",		-- colors: 47, 47, 47, 47
        440 => x"2F2F2F2F",		-- colors: 47, 47, 47, 47
        441 => x"2F2F2F2F",		-- colors: 47, 47, 47, 47
        442 => x"2F2F2F2F",		-- colors: 47, 47, 47, 47
        443 => x"2F2F2F2F",		-- colors: 47, 47, 47, 47
        444 => x"2F2F2F2F",		-- colors: 47, 47, 47, 47
        445 => x"2F2F2F2F",		-- colors: 47, 47, 47, 47
        446 => x"2F2F2F2F",		-- colors: 47, 47, 47, 47



--blue car sprite

                --  sprite 0
        447 => x"30303030",		-- colors: 48, 48, 48, 48
        448 => x"30303030",		-- colors: 48, 48, 48, 48
        449 => x"30303030",		-- colors: 48, 48, 48, 48
        450 => x"30303030",		-- colors: 48, 48, 48, 48
        451 => x"30303030",		-- colors: 48, 48, 48, 48
        452 => x"30303132",		-- colors: 48, 48, 49, 50
        453 => x"31303030",		-- colors: 49, 48, 48, 48
        454 => x"30303030",		-- colors: 48, 48, 48, 48
        455 => x"30303030",		-- colors: 48, 48, 48, 48
        456 => x"30303133",		-- colors: 48, 48, 49, 51
        457 => x"33333333",		-- colors: 51, 51, 51, 51
        458 => x"33333030",		-- colors: 51, 51, 48, 48
        459 => x"30303031",		-- colors: 48, 48, 48, 49
        460 => x"30303333",		-- colors: 48, 48, 51, 51
        461 => x"33333333",		-- colors: 51, 51, 51, 51
        462 => x"33333333",		-- colors: 51, 51, 51, 51
        463 => x"30303236",		-- colors: 48, 48, 50, 54
        464 => x"33333737",		-- colors: 51, 51, 55, 55
        465 => x"37373737",		-- colors: 55, 55, 55, 55
        466 => x"38383333",		-- colors: 56, 56, 51, 51
        467 => x"30303333",		-- colors: 48, 48, 51, 51
        468 => x"37373737",		-- colors: 55, 55, 55, 55
        469 => x"37373838",		-- colors: 55, 55, 56, 56
        470 => x"38383333",		-- colors: 56, 56, 51, 51
        471 => x"3C3C3737",		-- colors: 60, 60, 55, 55
        472 => x"37373737",		-- colors: 55, 55, 55, 55
        473 => x"38383838",		-- colors: 56, 56, 56, 56
        474 => x"38383333",		-- colors: 56, 56, 51, 51
        475 => x"33333737",		-- colors: 51, 51, 55, 55
        476 => x"37373738",		-- colors: 55, 55, 55, 56
        477 => x"38383838",		-- colors: 56, 56, 56, 56
        478 => x"38383333",		-- colors: 56, 56, 51, 51
        479 => x"33333737",		-- colors: 51, 51, 55, 55
        480 => x"37373738",		-- colors: 55, 55, 55, 56
        481 => x"38383838",		-- colors: 56, 56, 56, 56
        482 => x"38383333",		-- colors: 56, 56, 51, 51
        483 => x"33333737",		-- colors: 51, 51, 55, 55
        484 => x"37373744",		-- colors: 55, 55, 55, 68
        485 => x"38383838",		-- colors: 56, 56, 56, 56
        486 => x"38383333",		-- colors: 56, 56, 51, 51
        487 => x"3C3C3737",		-- colors: 60, 60, 55, 55
        488 => x"37373737",		-- colors: 55, 55, 55, 55
        489 => x"38383845",		-- colors: 56, 56, 56, 69
        490 => x"38383333",		-- colors: 56, 56, 51, 51
        491 => x"30303333",		-- colors: 48, 48, 51, 51
        492 => x"37373737",		-- colors: 55, 55, 55, 55
        493 => x"37373838",		-- colors: 55, 55, 56, 56
        494 => x"38383333",		-- colors: 56, 56, 51, 51
        495 => x"30313130",		-- colors: 48, 49, 49, 48
        496 => x"33333737",		-- colors: 51, 51, 55, 55
        497 => x"37373737",		-- colors: 55, 55, 55, 55
        498 => x"38383333",		-- colors: 56, 56, 51, 51
        499 => x"30303031",		-- colors: 48, 48, 48, 49
        500 => x"32483433",		-- colors: 50, 72, 52, 51
        501 => x"33333333",		-- colors: 51, 51, 51, 51
        502 => x"33333333",		-- colors: 51, 51, 51, 51
        503 => x"30303030",		-- colors: 48, 48, 48, 48
        504 => x"30303033",		-- colors: 48, 48, 48, 51
        505 => x"33333333",		-- colors: 51, 51, 51, 51
        506 => x"33333030",		-- colors: 51, 51, 48, 48
        507 => x"30303030",		-- colors: 48, 48, 48, 48
        508 => x"30303030",		-- colors: 48, 48, 48, 48
        509 => x"30303030",		-- colors: 48, 48, 48, 48
        510 => x"30303030",		-- colors: 48, 48, 48, 48

                --  sprite 1
        511 => x"30303030",		-- colors: 48, 48, 48, 48
        512 => x"30303030",		-- colors: 48, 48, 48, 48
        513 => x"30303030",		-- colors: 48, 48, 48, 48
        514 => x"30303030",		-- colors: 48, 48, 48, 48
        515 => x"30303030",		-- colors: 48, 48, 48, 48
        516 => x"30303232",		-- colors: 48, 48, 50, 50
        517 => x"31303030",		-- colors: 49, 48, 48, 48
        518 => x"30303030",		-- colors: 48, 48, 48, 48
        519 => x"30303031",		-- colors: 48, 48, 48, 49
        520 => x"30303333",		-- colors: 48, 48, 51, 51
        521 => x"30313130",		-- colors: 48, 49, 49, 48
        522 => x"30303030",		-- colors: 48, 48, 48, 48
        523 => x"34343533",		-- colors: 52, 52, 53, 51
        524 => x"33333333",		-- colors: 51, 51, 51, 51
        525 => x"33333031",		-- colors: 51, 51, 48, 49
        526 => x"32313030",		-- colors: 50, 49, 48, 48
        527 => x"37373333",		-- colors: 55, 55, 51, 51
        528 => x"37373737",		-- colors: 55, 55, 55, 55
        529 => x"33333933",		-- colors: 51, 51, 57, 51
        530 => x"333A3130",		-- colors: 51, 58, 49, 48
        531 => x"37373333",		-- colors: 55, 55, 51, 51
        532 => x"37373737",		-- colors: 55, 55, 55, 55
        533 => x"33333737",		-- colors: 51, 51, 55, 55
        534 => x"3B333331",		-- colors: 59, 51, 51, 49
        535 => x"33333333",		-- colors: 51, 51, 51, 51
        536 => x"3D3E3E3F",		-- colors: 61, 62, 62, 63
        537 => x"33333737",		-- colors: 51, 51, 55, 55
        538 => x"37373333",		-- colors: 55, 55, 51, 51
        539 => x"37373737",		-- colors: 55, 55, 55, 55
        540 => x"37373737",		-- colors: 55, 55, 55, 55
        541 => x"33333737",		-- colors: 51, 51, 55, 55
        542 => x"37373333",		-- colors: 55, 55, 51, 51
        543 => x"33404142",		-- colors: 51, 64, 65, 66
        544 => x"43373737",		-- colors: 67, 55, 55, 55
        545 => x"33333737",		-- colors: 51, 51, 55, 55
        546 => x"37373333",		-- colors: 55, 55, 51, 51
        547 => x"37373737",		-- colors: 55, 55, 55, 55
        548 => x"37373737",		-- colors: 55, 55, 55, 55
        549 => x"33333737",		-- colors: 51, 51, 55, 55
        550 => x"37373333",		-- colors: 55, 55, 51, 51
        551 => x"33333333",		-- colors: 51, 51, 51, 51
        552 => x"33333333",		-- colors: 51, 51, 51, 51
        553 => x"33333737",		-- colors: 51, 51, 55, 55
        554 => x"37373333",		-- colors: 55, 55, 51, 51
        555 => x"37373333",		-- colors: 55, 55, 51, 51
        556 => x"37373737",		-- colors: 55, 55, 55, 55
        557 => x"33333737",		-- colors: 51, 51, 55, 55
        558 => x"37334631",		-- colors: 55, 51, 70, 49
        559 => x"37373333",		-- colors: 55, 55, 51, 51
        560 => x"37373737",		-- colors: 55, 55, 55, 55
        561 => x"33473333",		-- colors: 51, 71, 51, 51
        562 => x"33333030",		-- colors: 51, 51, 48, 48
        563 => x"494A3530",		-- colors: 73, 74, 53, 48
        564 => x"33333333",		-- colors: 51, 51, 51, 51
        565 => x"33333030",		-- colors: 51, 51, 48, 48
        566 => x"31303030",		-- colors: 49, 48, 48, 48
        567 => x"30303031",		-- colors: 48, 48, 48, 49
        568 => x"31303333",		-- colors: 49, 48, 51, 51
        569 => x"33304B30",		-- colors: 51, 48, 75, 48
        570 => x"30303030",		-- colors: 48, 48, 48, 48
        571 => x"30303030",		-- colors: 48, 48, 48, 48
        572 => x"30313232",		-- colors: 48, 49, 50, 50
        573 => x"32313030",		-- colors: 50, 49, 48, 48
        574 => x"30303030",		-- colors: 48, 48, 48, 48
        
        
        
--red_car





       

--		****  MAP  ****
     
                --  sprite 0
        6992 => x"23232323",		-- colors: 35, 35, 35, 35
        6993 => x"23232323",		-- colors: 35, 35, 35, 35
        6994 => x"23232323",		-- colors: 35, 35, 35, 35
        6995 => x"23232323",		-- colors: 35, 35, 35, 35
        6996 => x"23232323",		-- colors: 35, 35, 35, 35
        6997 => x"23232323",		-- colors: 35, 35, 35, 35
        6998 => x"23232323",		-- colors: 35, 35, 35, 35
        6999 => x"23232323",		-- colors: 35, 35, 35, 35
        7000 => x"23232323",		-- colors: 35, 35, 35, 35
        7001 => x"23232323",		-- colors: 35, 35, 35, 35
        7002 => x"23232323",		-- colors: 35, 35, 35, 35
        7003 => x"23232323",		-- colors: 35, 35, 35, 35
        7004 => x"23232323",		-- colors: 35, 35, 35, 35
        7005 => x"23232323",		-- colors: 35, 35, 35, 35
        7006 => x"23232323",		-- colors: 35, 35, 35, 35
        7007 => x"23232323",		-- colors: 35, 35, 35, 35
        7008 => x"23232323",		-- colors: 35, 35, 35, 35
        7009 => x"23232323",		-- colors: 35, 35, 35, 35
        7010 => x"23232323",		-- colors: 35, 35, 35, 35
        7011 => x"23232323",		-- colors: 35, 35, 35, 35
        7012 => x"23232323",		-- colors: 35, 35, 35, 35
        7013 => x"23232323",		-- colors: 35, 35, 35, 35
        7014 => x"23232323",		-- colors: 35, 35, 35, 35
        7015 => x"23232323",		-- colors: 35, 35, 35, 35
        7016 => x"23232323",		-- colors: 35, 35, 35, 35
        7017 => x"23232323",		-- colors: 35, 35, 35, 35
        7018 => x"23232323",		-- colors: 35, 35, 35, 35
        7019 => x"23232323",		-- colors: 35, 35, 35, 35
        7020 => x"23232323",		-- colors: 35, 35, 35, 35
        7021 => x"23232323",		-- colors: 35, 35, 35, 35
        7022 => x"23232323",		-- colors: 35, 35, 35, 35
        7023 => x"23232323",		-- colors: 35, 35, 35, 35
        7024 => x"23232323",		-- colors: 35, 35, 35, 35
        7025 => x"23232323",		-- colors: 35, 35, 35, 35
        7026 => x"23232323",		-- colors: 35, 35, 35, 35
        7027 => x"23232323",		-- colors: 35, 35, 35, 35
        7028 => x"23232323",		-- colors: 35, 35, 35, 35
        7029 => x"23232323",		-- colors: 35, 35, 35, 35
        7030 => x"23232323",		-- colors: 35, 35, 35, 35
        7031 => x"23232323",		-- colors: 35, 35, 35, 35
        7032 => x"23232323",		-- colors: 35, 35, 35, 35
        7033 => x"23232323",		-- colors: 35, 35, 35, 35
        7034 => x"23232323",		-- colors: 35, 35, 35, 35
        7035 => x"23232323",		-- colors: 35, 35, 35, 35
        7036 => x"23232323",		-- colors: 35, 35, 35, 35
        7037 => x"23232323",		-- colors: 35, 35, 35, 35
        7038 => x"23232323",		-- colors: 35, 35, 35, 35
        7039 => x"23232323",		-- colors: 35, 35, 35, 35
        7040 => x"23232323",		-- colors: 35, 35, 35, 35
        7041 => x"23232323",		-- colors: 35, 35, 35, 35
        7042 => x"23232323",		-- colors: 35, 35, 35, 35
        7043 => x"23232323",		-- colors: 35, 35, 35, 35
        7044 => x"23232323",		-- colors: 35, 35, 35, 35
        7045 => x"23232323",		-- colors: 35, 35, 35, 35
        7046 => x"23232323",		-- colors: 35, 35, 35, 35
        7047 => x"23232323",		-- colors: 35, 35, 35, 35
        7048 => x"23232323",		-- colors: 35, 35, 35, 35
        7049 => x"23232323",		-- colors: 35, 35, 35, 35
        7050 => x"23232323",		-- colors: 35, 35, 35, 35
        7051 => x"23232323",		-- colors: 35, 35, 35, 35
        7052 => x"23232323",		-- colors: 35, 35, 35, 35
        7053 => x"23232323",		-- colors: 35, 35, 35, 35
        7054 => x"23232323",		-- colors: 35, 35, 35, 35
        7055 => x"23232323",		-- colors: 35, 35, 35, 35

                --  sprite 1
        7056 => x"24242424",		-- colors: 36, 36, 36, 36
        7057 => x"24242424",		-- colors: 36, 36, 36, 36
        7058 => x"24242424",		-- colors: 36, 36, 36, 36
        7059 => x"24242424",		-- colors: 36, 36, 36, 36
        7060 => x"24242424",		-- colors: 36, 36, 36, 36
        7061 => x"24242424",		-- colors: 36, 36, 36, 36
        7062 => x"24242424",		-- colors: 36, 36, 36, 36
        7063 => x"24242424",		-- colors: 36, 36, 36, 36
        7064 => x"24242424",		-- colors: 36, 36, 36, 36
        7065 => x"24242424",		-- colors: 36, 36, 36, 36
        7066 => x"24242424",		-- colors: 36, 36, 36, 36
        7067 => x"24242424",		-- colors: 36, 36, 36, 36
        7068 => x"24242424",		-- colors: 36, 36, 36, 36
        7069 => x"24242424",		-- colors: 36, 36, 36, 36
        7070 => x"24242424",		-- colors: 36, 36, 36, 36
        7071 => x"24242424",		-- colors: 36, 36, 36, 36
        7072 => x"24242424",		-- colors: 36, 36, 36, 36
        7073 => x"24242424",		-- colors: 36, 36, 36, 36
        7074 => x"24242424",		-- colors: 36, 36, 36, 36
        7075 => x"24242424",		-- colors: 36, 36, 36, 36
        7076 => x"24242424",		-- colors: 36, 36, 36, 36
        7077 => x"24242424",		-- colors: 36, 36, 36, 36
        7078 => x"24242424",		-- colors: 36, 36, 36, 36
        7079 => x"24242424",		-- colors: 36, 36, 36, 36
        7080 => x"24242424",		-- colors: 36, 36, 36, 36
        7081 => x"24242424",		-- colors: 36, 36, 36, 36
        7082 => x"24242424",		-- colors: 36, 36, 36, 36
        7083 => x"24242424",		-- colors: 36, 36, 36, 36
        7084 => x"24242424",		-- colors: 36, 36, 36, 36
        7085 => x"24242424",		-- colors: 36, 36, 36, 36
        7086 => x"24242424",		-- colors: 36, 36, 36, 36
        7087 => x"24242424",		-- colors: 36, 36, 36, 36
        7088 => x"24242424",		-- colors: 36, 36, 36, 36
        7089 => x"24242424",		-- colors: 36, 36, 36, 36
        7090 => x"24242424",		-- colors: 36, 36, 36, 36
        7091 => x"24242424",		-- colors: 36, 36, 36, 36
        7092 => x"24242424",		-- colors: 36, 36, 36, 36
        7093 => x"24242424",		-- colors: 36, 36, 36, 36
        7094 => x"24242424",		-- colors: 36, 36, 36, 36
        7095 => x"24242424",		-- colors: 36, 36, 36, 36
        7096 => x"24242424",		-- colors: 36, 36, 36, 36
        7097 => x"24242424",		-- colors: 36, 36, 36, 36
        7098 => x"24242424",		-- colors: 36, 36, 36, 36
        7099 => x"24242424",		-- colors: 36, 36, 36, 36
        7100 => x"24242424",		-- colors: 36, 36, 36, 36
        7101 => x"24242424",		-- colors: 36, 36, 36, 36
        7102 => x"24242424",		-- colors: 36, 36, 36, 36
        7103 => x"24242424",		-- colors: 36, 36, 36, 36
        7104 => x"24242424",		-- colors: 36, 36, 36, 36
        7105 => x"24242424",		-- colors: 36, 36, 36, 36
        7106 => x"24242424",		-- colors: 36, 36, 36, 36
        7107 => x"24242424",		-- colors: 36, 36, 36, 36
        7108 => x"24242424",		-- colors: 36, 36, 36, 36
        7109 => x"24242424",		-- colors: 36, 36, 36, 36
        7110 => x"24242424",		-- colors: 36, 36, 36, 36
        7111 => x"24242424",		-- colors: 36, 36, 36, 36
        7112 => x"24242424",		-- colors: 36, 36, 36, 36
        7113 => x"24242424",		-- colors: 36, 36, 36, 36
        7114 => x"24242424",		-- colors: 36, 36, 36, 36
        7115 => x"24242424",		-- colors: 36, 36, 36, 36
        7116 => x"24242424",		-- colors: 36, 36, 36, 36
        7117 => x"24242424",		-- colors: 36, 36, 36, 36
        7118 => x"24242424",		-- colors: 36, 36, 36, 36
        7119 => x"24242424",		-- colors: 36, 36, 36, 36

                --  sprite 2
        7120 => x"25252525",		-- colors: 37, 37, 37, 37
        7121 => x"25252525",		-- colors: 37, 37, 37, 37
        7122 => x"25252525",		-- colors: 37, 37, 37, 37
        7123 => x"25252525",		-- colors: 37, 37, 37, 37
        7124 => x"25252525",		-- colors: 37, 37, 37, 37
        7125 => x"25252525",		-- colors: 37, 37, 37, 37
        7126 => x"25252525",		-- colors: 37, 37, 37, 37
        7127 => x"25252525",		-- colors: 37, 37, 37, 37
        7128 => x"25252525",		-- colors: 37, 37, 37, 37
        7129 => x"25252525",		-- colors: 37, 37, 37, 37
        7130 => x"25252525",		-- colors: 37, 37, 37, 37
        7131 => x"25252525",		-- colors: 37, 37, 37, 37
        7132 => x"25252525",		-- colors: 37, 37, 37, 37
        7133 => x"25252525",		-- colors: 37, 37, 37, 37
        7134 => x"25252525",		-- colors: 37, 37, 37, 37
        7135 => x"25252525",		-- colors: 37, 37, 37, 37
        7136 => x"25252525",		-- colors: 37, 37, 37, 37
        7137 => x"25252525",		-- colors: 37, 37, 37, 37
        7138 => x"25252525",		-- colors: 37, 37, 37, 37
        7139 => x"25252525",		-- colors: 37, 37, 37, 37
        7140 => x"25252525",		-- colors: 37, 37, 37, 37
        7141 => x"25252525",		-- colors: 37, 37, 37, 37
        7142 => x"25252525",		-- colors: 37, 37, 37, 37
        7143 => x"25252525",		-- colors: 37, 37, 37, 37
        7144 => x"25252525",		-- colors: 37, 37, 37, 37
        7145 => x"25252525",		-- colors: 37, 37, 37, 37
        7146 => x"25252525",		-- colors: 37, 37, 37, 37
        7147 => x"25252525",		-- colors: 37, 37, 37, 37
        7148 => x"25252525",		-- colors: 37, 37, 37, 37
        7149 => x"25252525",		-- colors: 37, 37, 37, 37
        7150 => x"25252525",		-- colors: 37, 37, 37, 37
        7151 => x"25252525",		-- colors: 37, 37, 37, 37
        7152 => x"25252525",		-- colors: 37, 37, 37, 37
        7153 => x"25252525",		-- colors: 37, 37, 37, 37
        7154 => x"25252525",		-- colors: 37, 37, 37, 37
        7155 => x"25252525",		-- colors: 37, 37, 37, 37
        7156 => x"25252525",		-- colors: 37, 37, 37, 37
        7157 => x"25252525",		-- colors: 37, 37, 37, 37
        7158 => x"25252525",		-- colors: 37, 37, 37, 37
        7159 => x"25252525",		-- colors: 37, 37, 37, 37
        7160 => x"25252525",		-- colors: 37, 37, 37, 37
        7161 => x"25252525",		-- colors: 37, 37, 37, 37
        7162 => x"25252525",		-- colors: 37, 37, 37, 37
        7163 => x"25252525",		-- colors: 37, 37, 37, 37
        7164 => x"25252525",		-- colors: 37, 37, 37, 37
        7165 => x"25252525",		-- colors: 37, 37, 37, 37
        7166 => x"25252525",		-- colors: 37, 37, 37, 37
        7167 => x"25252525",		-- colors: 37, 37, 37, 37
        7168 => x"25252525",		-- colors: 37, 37, 37, 37
        7169 => x"25252525",		-- colors: 37, 37, 37, 37
        7170 => x"25252525",		-- colors: 37, 37, 37, 37
        7171 => x"25252525",		-- colors: 37, 37, 37, 37
        7172 => x"25252525",		-- colors: 37, 37, 37, 37
        7173 => x"25252525",		-- colors: 37, 37, 37, 37
        7174 => x"25252525",		-- colors: 37, 37, 37, 37
        7175 => x"25252525",		-- colors: 37, 37, 37, 37
        7176 => x"25252525",		-- colors: 37, 37, 37, 37
        7177 => x"25252525",		-- colors: 37, 37, 37, 37
        7178 => x"25252525",		-- colors: 37, 37, 37, 37
        7179 => x"25252525",		-- colors: 37, 37, 37, 37
        7180 => x"25252525",		-- colors: 37, 37, 37, 37
        7181 => x"25252525",		-- colors: 37, 37, 37, 37
        7182 => x"25252525",		-- colors: 37, 37, 37, 37
        7183 => x"25252525",		-- colors: 37, 37, 37, 37

                --  sprite 3
        7184 => x"26262626",		-- colors: 38, 38, 38, 38
        7185 => x"26262626",		-- colors: 38, 38, 38, 38
        7186 => x"26262626",		-- colors: 38, 38, 38, 38
        7187 => x"26262626",		-- colors: 38, 38, 38, 38
        7188 => x"26262626",		-- colors: 38, 38, 38, 38
        7189 => x"26262626",		-- colors: 38, 38, 38, 38
        7190 => x"26262626",		-- colors: 38, 38, 38, 38
        7191 => x"26262626",		-- colors: 38, 38, 38, 38
        7192 => x"26262626",		-- colors: 38, 38, 38, 38
        7193 => x"26262626",		-- colors: 38, 38, 38, 38
        7194 => x"26262626",		-- colors: 38, 38, 38, 38
        7195 => x"26262626",		-- colors: 38, 38, 38, 38
        7196 => x"26262626",		-- colors: 38, 38, 38, 38
        7197 => x"26262626",		-- colors: 38, 38, 38, 38
        7198 => x"26262626",		-- colors: 38, 38, 38, 38
        7199 => x"26262626",		-- colors: 38, 38, 38, 38
        7200 => x"26262626",		-- colors: 38, 38, 38, 38
        7201 => x"26262626",		-- colors: 38, 38, 38, 38
        7202 => x"26262626",		-- colors: 38, 38, 38, 38
        7203 => x"26262626",		-- colors: 38, 38, 38, 38
        7204 => x"26262626",		-- colors: 38, 38, 38, 38
        7205 => x"26262626",		-- colors: 38, 38, 38, 38
        7206 => x"26262626",		-- colors: 38, 38, 38, 38
        7207 => x"26262626",		-- colors: 38, 38, 38, 38
        7208 => x"26262626",		-- colors: 38, 38, 38, 38
        7209 => x"26262626",		-- colors: 38, 38, 38, 38
        7210 => x"26262626",		-- colors: 38, 38, 38, 38
        7211 => x"26262626",		-- colors: 38, 38, 38, 38
        7212 => x"26262626",		-- colors: 38, 38, 38, 38
        7213 => x"26262626",		-- colors: 38, 38, 38, 38
        7214 => x"26262626",		-- colors: 38, 38, 38, 38
        7215 => x"26262626",		-- colors: 38, 38, 38, 38
        7216 => x"26262626",		-- colors: 38, 38, 38, 38
        7217 => x"26262626",		-- colors: 38, 38, 38, 38
        7218 => x"26262626",		-- colors: 38, 38, 38, 38
        7219 => x"26262626",		-- colors: 38, 38, 38, 38
        7220 => x"26262626",		-- colors: 38, 38, 38, 38
        7221 => x"26262626",		-- colors: 38, 38, 38, 38
        7222 => x"26262626",		-- colors: 38, 38, 38, 38
        7223 => x"26262626",		-- colors: 38, 38, 38, 38
        7224 => x"26262626",		-- colors: 38, 38, 38, 38
        7225 => x"26262626",		-- colors: 38, 38, 38, 38
        7226 => x"26262626",		-- colors: 38, 38, 38, 38
        7227 => x"26262626",		-- colors: 38, 38, 38, 38
        7228 => x"26262626",		-- colors: 38, 38, 38, 38
        7229 => x"26262626",		-- colors: 38, 38, 38, 38
        7230 => x"26262626",		-- colors: 38, 38, 38, 38
        7231 => x"26262626",		-- colors: 38, 38, 38, 38
        7232 => x"26262626",		-- colors: 38, 38, 38, 38
        7233 => x"26262626",		-- colors: 38, 38, 38, 38
        7234 => x"26262626",		-- colors: 38, 38, 38, 38
        7235 => x"26262626",		-- colors: 38, 38, 38, 38
        7236 => x"26262626",		-- colors: 38, 38, 38, 38
        7237 => x"26262626",		-- colors: 38, 38, 38, 38
        7238 => x"26262626",		-- colors: 38, 38, 38, 38
        7239 => x"26262626",		-- colors: 38, 38, 38, 38
        7240 => x"26262626",		-- colors: 38, 38, 38, 38
        7241 => x"26262626",		-- colors: 38, 38, 38, 38
        7242 => x"26262626",		-- colors: 38, 38, 38, 38
        7243 => x"26262626",		-- colors: 38, 38, 38, 38
        7244 => x"26262626",		-- colors: 38, 38, 38, 38
        7245 => x"26262626",		-- colors: 38, 38, 38, 38
        7246 => x"26262626",		-- colors: 38, 38, 38, 38
        7247 => x"26262626",		-- colors: 38, 38, 38, 38

                --  sprite 4
        7248 => x"27272727",		-- colors: 39, 39, 39, 39
        7249 => x"27272827",		-- colors: 39, 39, 40, 39
        7250 => x"28292727",		-- colors: 40, 41, 39, 39
        7251 => x"27272727",		-- colors: 39, 39, 39, 39
        7252 => x"27272728",		-- colors: 39, 39, 39, 40
        7253 => x"28282828",		-- colors: 40, 40, 40, 40
        7254 => x"28282828",		-- colors: 40, 40, 40, 40
        7255 => x"27272727",		-- colors: 39, 39, 39, 39
        7256 => x"27272828",		-- colors: 39, 39, 40, 40
        7257 => x"28282A28",		-- colors: 40, 40, 42, 40
        7258 => x"28282828",		-- colors: 40, 40, 40, 40
        7259 => x"28272727",		-- colors: 40, 39, 39, 39
        7260 => x"27272828",		-- colors: 39, 39, 40, 40
        7261 => x"28282828",		-- colors: 40, 40, 40, 40
        7262 => x"2828282B",		-- colors: 40, 40, 40, 43
        7263 => x"28282727",		-- colors: 40, 40, 39, 39
        7264 => x"27272728",		-- colors: 39, 39, 39, 40
        7265 => x"28282828",		-- colors: 40, 40, 40, 40
        7266 => x"28282828",		-- colors: 40, 40, 40, 40
        7267 => x"28282827",		-- colors: 40, 40, 40, 39
        7268 => x"27272828",		-- colors: 39, 39, 40, 40
        7269 => x"28282828",		-- colors: 40, 40, 40, 40
        7270 => x"28282828",		-- colors: 40, 40, 40, 40
        7271 => x"28282827",		-- colors: 40, 40, 40, 39
        7272 => x"27282828",		-- colors: 39, 40, 40, 40
        7273 => x"28282828",		-- colors: 40, 40, 40, 40
        7274 => x"28282828",		-- colors: 40, 40, 40, 40
        7275 => x"28282727",		-- colors: 40, 40, 39, 39
        7276 => x"27282828",		-- colors: 39, 40, 40, 40
        7277 => x"28282828",		-- colors: 40, 40, 40, 40
        7278 => x"282C2828",		-- colors: 40, 44, 40, 40
        7279 => x"28282727",		-- colors: 40, 40, 39, 39
        7280 => x"27282828",		-- colors: 39, 40, 40, 40
        7281 => x"28282A2D",		-- colors: 40, 40, 42, 45
        7282 => x"2D282828",		-- colors: 45, 40, 40, 40
        7283 => x"28282727",		-- colors: 40, 40, 39, 39
        7284 => x"27272828",		-- colors: 39, 39, 40, 40
        7285 => x"282A282D",		-- colors: 40, 42, 40, 45
        7286 => x"2D282828",		-- colors: 45, 40, 40, 40
        7287 => x"28282727",		-- colors: 40, 40, 39, 39
        7288 => x"27272828",		-- colors: 39, 39, 40, 40
        7289 => x"28282828",		-- colors: 40, 40, 40, 40
        7290 => x"28282828",		-- colors: 40, 40, 40, 40
        7291 => x"27272727",		-- colors: 39, 39, 39, 39
        7292 => x"27272828",		-- colors: 39, 39, 40, 40
        7293 => x"28282828",		-- colors: 40, 40, 40, 40
        7294 => x"28282827",		-- colors: 40, 40, 40, 39
        7295 => x"27272727",		-- colors: 39, 39, 39, 39
        7296 => x"27272828",		-- colors: 39, 39, 40, 40
        7297 => x"28282828",		-- colors: 40, 40, 40, 40
        7298 => x"28282827",		-- colors: 40, 40, 40, 39
        7299 => x"27272727",		-- colors: 39, 39, 39, 39
        7300 => x"27272728",		-- colors: 39, 39, 39, 40
        7301 => x"27272828",		-- colors: 39, 39, 40, 40
        7302 => x"28282727",		-- colors: 40, 40, 39, 39
        7303 => x"27272727",		-- colors: 39, 39, 39, 39
        7304 => x"27272727",		-- colors: 39, 39, 39, 39
        7305 => x"27272828",		-- colors: 39, 39, 40, 40
        7306 => x"28272727",		-- colors: 40, 39, 39, 39
        7307 => x"27272727",		-- colors: 39, 39, 39, 39
        7308 => x"27272727",		-- colors: 39, 39, 39, 39
        7309 => x"27272727",		-- colors: 39, 39, 39, 39
        7310 => x"27272727",		-- colors: 39, 39, 39, 39
        7311 => x"27272727",		-- colors: 39, 39, 39, 39
others => x"00000000"
	);


begin

	process(i_clk)
	begin
		if rising_edge(i_clk) then
			-- memory write --
			if i_we = '1' then
				mem(to_integer(unsigned(i_w_addr))) <= i_data;
			end if;
			-- memory read -- 
			o_data <= mem(to_integer(unsigned(i_r_addr)));
			
		end if; 
	end process;

end architecture arch;
