
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity ram is
	generic
	(
		DATA_WIDTH : natural := 32;		    -- 4 byte one line of memory
		ADDR_WIDTH : natural := 13			    -- 24576 bytes size of memory
	);

	port(
		i_clk    : in  std_logic;
		i_r_addr : in  std_logic_vector(ADDR_WIDTH-1 downto 0);
		i_data   : in  std_logic_vector(DATA_WIDTH-1 downto 0);
		i_we     : in  std_logic;
		i_w_addr : in  std_logic_vector(ADDR_WIDTH-1 downto 0);
		o_data   : out std_logic_vector(DATA_WIDTH-1 downto 0)
	);
end entity ram;

architecture arch of ram is

	type ram_t is array (0 to 2**ADDR_WIDTH-1) of std_logic_vector(DATA_WIDTH-1 downto 0);


-- GENERATED BY BC_MEM_PACKER

-- DATE: Thu May 18 16:01:02 2017

	signal mem : ram_t := (

--			***** COLOR PALLETE *****


--kirby colors

			0 => x"00000000",
			1 => x"00ea8bff",
			2 => x"00e98afe",
			3 => x"003d3d40",
			4 => x"00811699",
			5 => x"00ea8aff",
			6 => x"000303d5",

--mapa colors

			7 => x"00353b39",
			8 => x"000bac82",
			9 => x"00000000",
			10 => x"0018704c",
			11 => x"000aab81",
			12 => x"000cac83",
			13 => x"000cad83",
			14 => x"000cac82",
			15 => x"00ffffff",
	

--red_car

			16 => x"00353b39",
			17 => x"0007072c",
			18 => x"000000fe",
			19 => x"0008072c",
			20 => x"00b19357",
			21 => x"000800fe",
			22 => x"0000dcd6",
			23 => x"0012082c",
			24 => x"0019092c",
			25 => x"0016092c",
			26 => x"001d01fb",

--blue_car
                
      27 => x"00353b39",
		28 => x"0008072c",
		29 => x"00ab1c2b",
		30 => x"00b09256",
		31 => x"0000dcd6",
		32 => x"000e082c",
  
                
					 
--			***** 16x16 IMAGES *****
--			OVERWORLD SPRITES
        
--kirby sprites        
               
--  sprite 0

        255 => x"00000000",		-- colors: 0, 0, 0, 0
        256 => x"00000000",		-- colors: 0, 0, 0, 0
        257 => x"00000000",		-- colors: 0, 0, 0, 0
        258 => x"00000000",		-- colors: 0, 0, 0, 0
        259 => x"00000000",		-- colors: 0, 0, 0, 0
        260 => x"00000000",		-- colors: 0, 0, 0, 0
        261 => x"00000000",		-- colors: 0, 0, 0, 0
        262 => x"00000000",		-- colors: 0, 0, 0, 0
        263 => x"00000000",		-- colors: 0, 0, 0, 0
        264 => x"00000000",		-- colors: 0, 0, 0, 0
        265 => x"00000000",		-- colors: 0, 0, 0, 0
        266 => x"00000000",		-- colors: 0, 0, 0, 0
        267 => x"00000000",		-- colors: 0, 0, 0, 0
        268 => x"00000000",		-- colors: 0, 0, 0, 0
        269 => x"00000000",		-- colors: 0, 0, 0, 0
        270 => x"00000000",		-- colors: 0, 0, 0, 0
        271 => x"00000000",		-- colors: 0, 0, 0, 0
        272 => x"00000000",		-- colors: 0, 0, 0, 0
        273 => x"00000000",		-- colors: 0, 0, 0, 0
        274 => x"00000000",		-- colors: 0, 0, 0, 0
        275 => x"00000000",		-- colors: 0, 0, 0, 0
        276 => x"00000000",		-- colors: 0, 0, 0, 0
        277 => x"00000000",		-- colors: 0, 0, 0, 0
        278 => x"00000000",		-- colors: 0, 0, 0, 0
        279 => x"00000000",		-- colors: 0, 0, 0, 0
        280 => x"00000000",		-- colors: 0, 0, 0, 0
        281 => x"00000000",		-- colors: 0, 0, 0, 0
        282 => x"00000000",		-- colors: 0, 0, 0, 0
        283 => x"00000000",		-- colors: 0, 0, 0, 0
        284 => x"00000101",		-- colors: 0, 0, 1, 1
        285 => x"01020000",		-- colors: 1, 2, 0, 0
        286 => x"00000000",		-- colors: 0, 0, 0, 0
        287 => x"00000000",		-- colors: 0, 0, 0, 0
        288 => x"00010101",		-- colors: 0, 1, 1, 1
        289 => x"01010100",		-- colors: 1, 1, 1, 0
        290 => x"00000000",		-- colors: 0, 0, 0, 0
        291 => x"00000000",		-- colors: 0, 0, 0, 0
        292 => x"01010301",		-- colors: 1, 1, 3, 1
        293 => x"01030101",		-- colors: 1, 3, 1, 1
        294 => x"00000000",		-- colors: 0, 0, 0, 0
        295 => x"00000001",		-- colors: 0, 0, 0, 1
        296 => x"01010301",		-- colors: 1, 1, 3, 1
        297 => x"01030101",		-- colors: 1, 3, 1, 1
        298 => x"01000000",		-- colors: 1, 0, 0, 0
        299 => x"00000001",		-- colors: 0, 0, 0, 1
        300 => x"01040101",		-- colors: 1, 4, 1, 1
        301 => x"01010401",		-- colors: 1, 1, 4, 1
        302 => x"01000000",		-- colors: 1, 0, 0, 0
        303 => x"00000000",		-- colors: 0, 0, 0, 0
        304 => x"05010101",		-- colors: 5, 1, 1, 1
        305 => x"01010101",		-- colors: 1, 1, 1, 1
        306 => x"00000000",		-- colors: 0, 0, 0, 0
        307 => x"00000000",		-- colors: 0, 0, 0, 0
        308 => x"00010101",		-- colors: 0, 1, 1, 1
        309 => x"01010100",		-- colors: 1, 1, 1, 0
        310 => x"00000000",		-- colors: 0, 0, 0, 0
        311 => x"00000000",		-- colors: 0, 0, 0, 0
        312 => x"00000101",		-- colors: 0, 0, 1, 1
        313 => x"01010000",		-- colors: 1, 1, 0, 0
        314 => x"00000000",		-- colors: 0, 0, 0, 0
        315 => x"00000000",		-- colors: 0, 0, 0, 0
        316 => x"00060600",		-- colors: 0, 6, 6, 0
        317 => x"00060600",		-- colors: 0, 6, 6, 0
        318 => x"00000000",		-- colors: 0, 0, 0, 0
        

        
--red_car sprite



        
                --  sprite 0
        447 => x"10101010",		-- colors: 16, 16, 16, 16
        448 => x"10101010",		-- colors: 16, 16, 16, 16
        449 => x"10101010",		-- colors: 16, 16, 16, 16
        450 => x"10101010",		-- colors: 16, 16, 16, 16
        451 => x"10101010",		-- colors: 16, 16, 16, 16
        452 => x"10101111",		-- colors: 16, 16, 17, 17
        453 => x"11111110",		-- colors: 17, 17, 17, 16
        454 => x"10101010",		-- colors: 16, 16, 16, 16
        455 => x"10101010",		-- colors: 16, 16, 16, 16
        456 => x"10101111",		-- colors: 16, 16, 17, 17
        457 => x"11111111",		-- colors: 17, 17, 17, 17
        458 => x"10101010",		-- colors: 16, 16, 16, 16
        459 => x"10101111",		-- colors: 16, 16, 17, 17
        460 => x"11111111",		-- colors: 17, 17, 17, 17
        461 => x"12121212",		-- colors: 18, 18, 18, 18
        462 => x"13131212",		-- colors: 19, 19, 18, 18
        463 => x"10111112",		-- colors: 16, 17, 17, 18
        464 => x"12121111",		-- colors: 18, 18, 17, 17
        465 => x"12121212",		-- colors: 18, 18, 18, 18
        466 => x"13131212",		-- colors: 19, 19, 18, 18
        467 => x"11111512",		-- colors: 17, 17, 21, 18
        468 => x"12121111",		-- colors: 18, 18, 17, 17
        469 => x"13131313",		-- colors: 19, 19, 19, 19
        470 => x"13131313",		-- colors: 19, 19, 19, 19
        471 => x"11111212",		-- colors: 17, 17, 18, 18
        472 => x"12121111",		-- colors: 18, 18, 17, 17
        473 => x"12121212",		-- colors: 18, 18, 18, 18
        474 => x"12121212",		-- colors: 18, 18, 18, 18
        475 => x"11111212",		-- colors: 17, 17, 18, 18
        476 => x"12121111",		-- colors: 18, 18, 17, 17
        477 => x"12121212",		-- colors: 18, 18, 18, 18
        478 => x"12121213",		-- colors: 18, 18, 18, 19
        479 => x"11111212",		-- colors: 17, 17, 18, 18
        480 => x"12121111",		-- colors: 18, 18, 17, 17
        481 => x"12121212",		-- colors: 18, 18, 18, 18
        482 => x"12121212",		-- colors: 18, 18, 18, 18
        483 => x"11111212",		-- colors: 17, 17, 18, 18
        484 => x"12121111",		-- colors: 18, 18, 17, 17
        485 => x"17181819",		-- colors: 23, 24, 24, 25
        486 => x"13131313",		-- colors: 19, 19, 19, 19
        487 => x"10111112",		-- colors: 16, 17, 17, 18
        488 => x"12121111",		-- colors: 18, 18, 17, 17
        489 => x"12121212",		-- colors: 18, 18, 18, 18
        490 => x"13131212",		-- colors: 19, 19, 18, 18
        491 => x"10101111",		-- colors: 16, 16, 17, 17
        492 => x"11111111",		-- colors: 17, 17, 17, 17
        493 => x"12121212",		-- colors: 18, 18, 18, 18
        494 => x"13131212",		-- colors: 19, 19, 18, 18
        495 => x"10101010",		-- colors: 16, 16, 16, 16
        496 => x"10101111",		-- colors: 16, 16, 17, 17
        497 => x"11111111",		-- colors: 17, 17, 17, 17
        498 => x"10101010",		-- colors: 16, 16, 16, 16
        499 => x"10101010",		-- colors: 16, 16, 16, 16
        500 => x"10101111",		-- colors: 16, 16, 17, 17
        501 => x"11111110",		-- colors: 17, 17, 17, 16
        502 => x"10101010",		-- colors: 16, 16, 16, 16
        503 => x"10101010",		-- colors: 16, 16, 16, 16
        504 => x"10101010",		-- colors: 16, 16, 16, 16
        505 => x"10101010",		-- colors: 16, 16, 16, 16
        506 => x"10101010",		-- colors: 16, 16, 16, 16
        507 => x"10101010",		-- colors: 16, 16, 16, 16
        508 => x"10101010",		-- colors: 16, 16, 16, 16
        509 => x"10101010",		-- colors: 16, 16, 16, 16
        510 => x"10101010",		-- colors: 16, 16, 16, 16

                --  sprite 1
        511 => x"10101010",		-- colors: 16, 16, 16, 16
        512 => x"10101010",		-- colors: 16, 16, 16, 16
        513 => x"10101010",		-- colors: 16, 16, 16, 16
        514 => x"10101010",		-- colors: 16, 16, 16, 16
        515 => x"10101111",		-- colors: 16, 16, 17, 17
        516 => x"11111111",		-- colors: 17, 17, 17, 17
        517 => x"11101010",		-- colors: 17, 16, 16, 16
        518 => x"10101010",		-- colors: 16, 16, 16, 16
        519 => x"11111111",		-- colors: 17, 17, 17, 17
        520 => x"11111111",		-- colors: 17, 17, 17, 17
        521 => x"11111010",		-- colors: 17, 17, 16, 16
        522 => x"10101010",		-- colors: 16, 16, 16, 16
        523 => x"11111414",		-- colors: 17, 17, 20, 20
        524 => x"12121212",		-- colors: 18, 18, 18, 18
        525 => x"12121111",		-- colors: 18, 18, 17, 17
        526 => x"10101010",		-- colors: 16, 16, 16, 16
        527 => x"11111414",		-- colors: 17, 17, 20, 20
        528 => x"14141212",		-- colors: 20, 20, 18, 18
        529 => x"12121212",		-- colors: 18, 18, 18, 18
        530 => x"11111010",		-- colors: 17, 17, 16, 16
        531 => x"11111414",		-- colors: 17, 17, 20, 20
        532 => x"14141414",		-- colors: 20, 20, 20, 20
        533 => x"12121212",		-- colors: 18, 18, 18, 18
        534 => x"12121616",		-- colors: 18, 18, 22, 22
        535 => x"11111414",		-- colors: 17, 17, 20, 20
        536 => x"14141414",		-- colors: 20, 20, 20, 20
        537 => x"14121212",		-- colors: 20, 18, 18, 18
        538 => x"12121111",		-- colors: 18, 18, 17, 17
        539 => x"11111414",		-- colors: 17, 17, 20, 20
        540 => x"14141414",		-- colors: 20, 20, 20, 20
        541 => x"14121212",		-- colors: 20, 18, 18, 18
        542 => x"12121111",		-- colors: 18, 18, 17, 17
        543 => x"11111414",		-- colors: 17, 17, 20, 20
        544 => x"14141414",		-- colors: 20, 20, 20, 20
        545 => x"14121212",		-- colors: 20, 18, 18, 18
        546 => x"12121111",		-- colors: 18, 18, 17, 17
        547 => x"11111414",		-- colors: 17, 17, 20, 20
        548 => x"14141414",		-- colors: 20, 20, 20, 20
        549 => x"12121212",		-- colors: 18, 18, 18, 18
        550 => x"12121616",		-- colors: 18, 18, 22, 22
        551 => x"11111414",		-- colors: 17, 17, 20, 20
        552 => x"14141A12",		-- colors: 20, 20, 26, 18
        553 => x"12121212",		-- colors: 18, 18, 18, 18
        554 => x"11111010",		-- colors: 17, 17, 16, 16
        555 => x"11111414",		-- colors: 17, 17, 20, 20
        556 => x"12121212",		-- colors: 18, 18, 18, 18
        557 => x"12121111",		-- colors: 18, 18, 17, 17
        558 => x"10101010",		-- colors: 16, 16, 16, 16
        559 => x"11111111",		-- colors: 17, 17, 17, 17
        560 => x"11111111",		-- colors: 17, 17, 17, 17
        561 => x"11111010",		-- colors: 17, 17, 16, 16
        562 => x"10101010",		-- colors: 16, 16, 16, 16
        563 => x"10101111",		-- colors: 16, 16, 17, 17
        564 => x"11111111",		-- colors: 17, 17, 17, 17
        565 => x"11101010",		-- colors: 17, 16, 16, 16
        566 => x"10101010",		-- colors: 16, 16, 16, 16
        567 => x"10101010",		-- colors: 16, 16, 16, 16
        568 => x"10101010",		-- colors: 16, 16, 16, 16
        569 => x"10101010",		-- colors: 16, 16, 16, 16
        570 => x"10101010",		-- colors: 16, 16, 16, 16
        571 => x"10101010",		-- colors: 16, 16, 16, 16
        572 => x"10101010",		-- colors: 16, 16, 16, 16
        573 => x"10101010",		-- colors: 16, 16, 16, 16
        574 => x"10101010",		-- colors: 16, 16, 16, 16
--blue car sprite

       
                --  sprite 0
        575 => x"1B1B1B1B",		-- colors: 27, 27, 27, 27
        576 => x"1B1B1B1B",		-- colors: 27, 27, 27, 27
        577 => x"1B1B1B1B",		-- colors: 27, 27, 27, 27
        578 => x"1B1B1B1B",		-- colors: 27, 27, 27, 27
        579 => x"1B1B1B1B",		-- colors: 27, 27, 27, 27
        580 => x"1B1B1B1B",		-- colors: 27, 27, 27, 27
        581 => x"1B1B1B1B",		-- colors: 27, 27, 27, 27
        582 => x"1B1B1B1B",		-- colors: 27, 27, 27, 27
        583 => x"1B1B1B1B",		-- colors: 27, 27, 27, 27
        584 => x"1B1B1B1C",		-- colors: 27, 27, 27, 28
        585 => x"1C1C1C1C",		-- colors: 28, 28, 28, 28
        586 => x"1C1C1B1B",		-- colors: 28, 28, 27, 27
        587 => x"1B1B1B1B",		-- colors: 27, 27, 27, 27
        588 => x"1B1B1C1C",		-- colors: 27, 27, 28, 28
        589 => x"1C1C1C1C",		-- colors: 28, 28, 28, 28
        590 => x"1C1C1C1C",		-- colors: 28, 28, 28, 28
        591 => x"1B1B1B1B",		-- colors: 27, 27, 27, 27
        592 => x"1C1C1D1D",		-- colors: 28, 28, 29, 29
        593 => x"1D1D1D1D",		-- colors: 29, 29, 29, 29
        594 => x"1E1E1C1C",		-- colors: 30, 30, 28, 28
        595 => x"1B1B1C1C",		-- colors: 27, 27, 28, 28
        596 => x"1D1D1D1D",		-- colors: 29, 29, 29, 29
        597 => x"1D1D1E1E",		-- colors: 29, 29, 30, 30
        598 => x"1E1E1C1C",		-- colors: 30, 30, 28, 28
        599 => x"1F1F1D1D",		-- colors: 31, 31, 29, 29
        600 => x"1D1D1D1D",		-- colors: 29, 29, 29, 29
        601 => x"1E1E1E1E",		-- colors: 30, 30, 30, 30
        602 => x"1E1E1C1C",		-- colors: 30, 30, 28, 28
        603 => x"1C1C1D1D",		-- colors: 28, 28, 29, 29
        604 => x"1D1D1D1E",		-- colors: 29, 29, 29, 30
        605 => x"1E1E1E1E",		-- colors: 30, 30, 30, 30
        606 => x"1E1E1C1C",		-- colors: 30, 30, 28, 28
        607 => x"1C1C1D1D",		-- colors: 28, 28, 29, 29
        608 => x"1D1D1D1E",		-- colors: 29, 29, 29, 30
        609 => x"1E1E1E1E",		-- colors: 30, 30, 30, 30
        610 => x"1E1E1C1C",		-- colors: 30, 30, 28, 28
        611 => x"1C1C1D1D",		-- colors: 28, 28, 29, 29
        612 => x"1D1D1D1E",		-- colors: 29, 29, 29, 30
        613 => x"1E1E1E1E",		-- colors: 30, 30, 30, 30
        614 => x"1E1E1C1C",		-- colors: 30, 30, 28, 28
        615 => x"1F1F1D1D",		-- colors: 31, 31, 29, 29
        616 => x"1D1D1D1D",		-- colors: 29, 29, 29, 29
        617 => x"1E1E1E1E",		-- colors: 30, 30, 30, 30
        618 => x"1E1E1C1C",		-- colors: 30, 30, 28, 28
        619 => x"1B1B1C1C",		-- colors: 27, 27, 28, 28
        620 => x"1D1D1D1D",		-- colors: 29, 29, 29, 29
        621 => x"1D1D1E1E",		-- colors: 29, 29, 30, 30
        622 => x"1E1E1C1C",		-- colors: 30, 30, 28, 28
        623 => x"1B1B1B1B",		-- colors: 27, 27, 27, 27
        624 => x"1C1C1D1D",		-- colors: 28, 28, 29, 29
        625 => x"1D1D1D1D",		-- colors: 29, 29, 29, 29
        626 => x"1E1E1C1C",		-- colors: 30, 30, 28, 28
        627 => x"1B1B1B1B",		-- colors: 27, 27, 27, 27
        628 => x"1B1B1C1C",		-- colors: 27, 27, 28, 28
        629 => x"1C1C1C1C",		-- colors: 28, 28, 28, 28
        630 => x"1C1C1C1C",		-- colors: 28, 28, 28, 28
        631 => x"1B1B1B1B",		-- colors: 27, 27, 27, 27
        632 => x"1B1B1B1C",		-- colors: 27, 27, 27, 28
        633 => x"1C1C1C1C",		-- colors: 28, 28, 28, 28
        634 => x"1C1C1B1B",		-- colors: 28, 28, 27, 27
        635 => x"1B1B1B1B",		-- colors: 27, 27, 27, 27
        636 => x"1B1B1B1B",		-- colors: 27, 27, 27, 27
        637 => x"1B1B1B1B",		-- colors: 27, 27, 27, 27
        638 => x"1B1B1B1B",		-- colors: 27, 27, 27, 27

                --  sprite 1
        639 => x"1B1B1B1B",		-- colors: 27, 27, 27, 27
        640 => x"1B1B1B1B",		-- colors: 27, 27, 27, 27
        641 => x"1B1B1B1B",		-- colors: 27, 27, 27, 27
        642 => x"1B1B1B1B",		-- colors: 27, 27, 27, 27
        643 => x"1B1B1B1B",		-- colors: 27, 27, 27, 27
        644 => x"1B1B1B1B",		-- colors: 27, 27, 27, 27
        645 => x"1B1B1B1B",		-- colors: 27, 27, 27, 27
        646 => x"1B1B1B1B",		-- colors: 27, 27, 27, 27
        647 => x"1B1B1B1B",		-- colors: 27, 27, 27, 27
        648 => x"1B1B1C1C",		-- colors: 27, 27, 28, 28
        649 => x"1C1B1B1B",		-- colors: 28, 27, 27, 27
        650 => x"1B1B1B1B",		-- colors: 27, 27, 27, 27
        651 => x"1B1B1B1B",		-- colors: 27, 27, 27, 27
        652 => x"1C1C1C1C",		-- colors: 28, 28, 28, 28
        653 => x"1C1C1B1B",		-- colors: 28, 28, 27, 27
        654 => x"1B1B1B1B",		-- colors: 27, 27, 27, 27
        655 => x"1D1D1C1C",		-- colors: 29, 29, 28, 28
        656 => x"1D1D1D1D",		-- colors: 29, 29, 29, 29
        657 => x"1C1C1C1C",		-- colors: 28, 28, 28, 28
        658 => x"1C1C1B1B",		-- colors: 28, 28, 27, 27
        659 => x"1D1D1C1C",		-- colors: 29, 29, 28, 28
        660 => x"1D1D1D1D",		-- colors: 29, 29, 29, 29
        661 => x"1C1C1D1D",		-- colors: 28, 28, 29, 29
        662 => x"1D1C1C1B",		-- colors: 29, 28, 28, 27
        663 => x"1C1C1C1C",		-- colors: 28, 28, 28, 28
        664 => x"1C20201C",		-- colors: 28, 32, 32, 28
        665 => x"1C1C1D1D",		-- colors: 28, 28, 29, 29
        666 => x"1D1D1C1C",		-- colors: 29, 29, 28, 28
        667 => x"1D1D1D1D",		-- colors: 29, 29, 29, 29
        668 => x"1D1D1D1D",		-- colors: 29, 29, 29, 29
        669 => x"1C1C1D1D",		-- colors: 28, 28, 29, 29
        670 => x"1D1D1C1C",		-- colors: 29, 29, 28, 28
        671 => x"1C1D1D1D",		-- colors: 28, 29, 29, 29
        672 => x"1D1D1D1D",		-- colors: 29, 29, 29, 29
        673 => x"1C1C1D1D",		-- colors: 28, 28, 29, 29
        674 => x"1D1D1C1C",		-- colors: 29, 29, 28, 28
        675 => x"1D1D1D1D",		-- colors: 29, 29, 29, 29
        676 => x"1D1D1D1D",		-- colors: 29, 29, 29, 29
        677 => x"1C1C1D1D",		-- colors: 28, 28, 29, 29
        678 => x"1D1D1C1C",		-- colors: 29, 29, 28, 28
        679 => x"1C1C1C1C",		-- colors: 28, 28, 28, 28
        680 => x"1C1C1C1C",		-- colors: 28, 28, 28, 28
        681 => x"1C1C1D1D",		-- colors: 28, 28, 29, 29
        682 => x"1D1D1C1C",		-- colors: 29, 29, 28, 28
        683 => x"1D1D1C1C",		-- colors: 29, 29, 28, 28
        684 => x"1D1D1D1D",		-- colors: 29, 29, 29, 29
        685 => x"1C1C1D1D",		-- colors: 28, 28, 29, 29
        686 => x"1D1C1C1B",		-- colors: 29, 28, 28, 27
        687 => x"1D1D1C1C",		-- colors: 29, 29, 28, 28
        688 => x"1D1D1D1D",		-- colors: 29, 29, 29, 29
        689 => x"1C1C1C1C",		-- colors: 28, 28, 28, 28
        690 => x"1C1C1B1B",		-- colors: 28, 28, 27, 27
        691 => x"1B1B1B1B",		-- colors: 27, 27, 27, 27
        692 => x"1C1C1C1C",		-- colors: 28, 28, 28, 28
        693 => x"1C1C1B1B",		-- colors: 28, 28, 27, 27
        694 => x"1B1B1B1B",		-- colors: 27, 27, 27, 27
        695 => x"1B1B1B1B",		-- colors: 27, 27, 27, 27
        696 => x"1B1B1C1C",		-- colors: 27, 27, 28, 28
        697 => x"1C1B1B1B",		-- colors: 28, 27, 27, 27
        698 => x"1B1B1B1B",		-- colors: 27, 27, 27, 27
        699 => x"1B1B1B1B",		-- colors: 27, 27, 27, 27
        700 => x"1B1B1B1B",		-- colors: 27, 27, 27, 27
        701 => x"1B1B1B1B",		-- colors: 27, 27, 27, 27
        702 => x"1B1B1B1B",		-- colors: 27, 27, 27, 27
 
--		****  MAP  ****
            
        
                --  sprite 0
        1000 => x"07070707",		-- colors: 7, 7, 7, 7
        1001 => x"07070707",		-- colors: 7, 7, 7, 7
        1002 => x"07070707",		-- colors: 7, 7, 7, 7
        1003 => x"07070707",		-- colors: 7, 7, 7, 7
        1004 => x"07070707",		-- colors: 7, 7, 7, 7
        1005 => x"07070707",		-- colors: 7, 7, 7, 7
        1006 => x"07070707",		-- colors: 7, 7, 7, 7
        1007 => x"07070707",		-- colors: 7, 7, 7, 7
        1008 => x"07070707",		-- colors: 7, 7, 7, 7
        1009 => x"07070707",		-- colors: 7, 7, 7, 7
        1010 => x"07070707",		-- colors: 7, 7, 7, 7
        1011 => x"07070707",		-- colors: 7, 7, 7, 7
        1012 => x"07070707",		-- colors: 7, 7, 7, 7
        1013 => x"07070707",		-- colors: 7, 7, 7, 7
        1014 => x"07070707",		-- colors: 7, 7, 7, 7
        1015 => x"07070707",		-- colors: 7, 7, 7, 7
        1016 => x"07070707",		-- colors: 7, 7, 7, 7
        1017 => x"07070707",		-- colors: 7, 7, 7, 7
        1018 => x"07070707",		-- colors: 7, 7, 7, 7
        1019 => x"07070707",		-- colors: 7, 7, 7, 7
        1020 => x"07070707",		-- colors: 7, 7, 7, 7
        1021 => x"07070707",		-- colors: 7, 7, 7, 7
        1022 => x"07070707",		-- colors: 7, 7, 7, 7
        1023 => x"07070707",		-- colors: 7, 7, 7, 7
        1024 => x"07070707",		-- colors: 7, 7, 7, 7
        1025 => x"07070707",		-- colors: 7, 7, 7, 7
        1026 => x"07070707",		-- colors: 7, 7, 7, 7
        1027 => x"07070707",		-- colors: 7, 7, 7, 7
        1028 => x"07070707",		-- colors: 7, 7, 7, 7
        1029 => x"07070707",		-- colors: 7, 7, 7, 7
        1030 => x"07070707",		-- colors: 7, 7, 7, 7
        1031 => x"07070707",		-- colors: 7, 7, 7, 7
        1032 => x"07070707",		-- colors: 7, 7, 7, 7
        1033 => x"07070707",		-- colors: 7, 7, 7, 7
        1034 => x"07070707",		-- colors: 7, 7, 7, 7
        1035 => x"07070707",		-- colors: 7, 7, 7, 7
        1036 => x"07070707",		-- colors: 7, 7, 7, 7
        1037 => x"07070707",		-- colors: 7, 7, 7, 7
        1038 => x"07070707",		-- colors: 7, 7, 7, 7
        1039 => x"07070707",		-- colors: 7, 7, 7, 7
        1040 => x"07070707",		-- colors: 7, 7, 7, 7
        1041 => x"07070707",		-- colors: 7, 7, 7, 7
        1042 => x"07070707",		-- colors: 7, 7, 7, 7
        1043 => x"07070707",		-- colors: 7, 7, 7, 7
        1044 => x"07070707",		-- colors: 7, 7, 7, 7
        1045 => x"07070707",		-- colors: 7, 7, 7, 7
        1046 => x"07070707",		-- colors: 7, 7, 7, 7
        1047 => x"07070707",		-- colors: 7, 7, 7, 7
        1048 => x"07070707",		-- colors: 7, 7, 7, 7
        1049 => x"07070707",		-- colors: 7, 7, 7, 7
        1050 => x"07070707",		-- colors: 7, 7, 7, 7
        1051 => x"07070707",		-- colors: 7, 7, 7, 7
        1052 => x"07070707",		-- colors: 7, 7, 7, 7
        1053 => x"07070707",		-- colors: 7, 7, 7, 7
        1054 => x"07070707",		-- colors: 7, 7, 7, 7
        1055 => x"07070707",		-- colors: 7, 7, 7, 7
        1056 => x"07070707",		-- colors: 7, 7, 7, 7
        1057 => x"07070707",		-- colors: 7, 7, 7, 7
        1058 => x"07070707",		-- colors: 7, 7, 7, 7
        1059 => x"07070707",		-- colors: 7, 7, 7, 7
        1060 => x"07070707",		-- colors: 7, 7, 7, 7
        1061 => x"07070707",		-- colors: 7, 7, 7, 7
        1062 => x"07070707",		-- colors: 7, 7, 7, 7
        1063 => x"07070707",		-- colors: 7, 7, 7, 7

                --  sprite 1
        1064 => x"08080808",		-- colors: 8, 8, 8, 8
        1065 => x"08080808",		-- colors: 8, 8, 8, 8
        1066 => x"08080808",		-- colors: 8, 8, 8, 8
        1067 => x"08080808",		-- colors: 8, 8, 8, 8
        1068 => x"08080808",		-- colors: 8, 8, 8, 8
        1069 => x"08080808",		-- colors: 8, 8, 8, 8
        1070 => x"08080808",		-- colors: 8, 8, 8, 8
        1071 => x"08080808",		-- colors: 8, 8, 8, 8
        1072 => x"08080808",		-- colors: 8, 8, 8, 8
        1073 => x"08080808",		-- colors: 8, 8, 8, 8
        1074 => x"08080808",		-- colors: 8, 8, 8, 8
        1075 => x"08080808",		-- colors: 8, 8, 8, 8
        1076 => x"08080808",		-- colors: 8, 8, 8, 8
        1077 => x"08080808",		-- colors: 8, 8, 8, 8
        1078 => x"08080808",		-- colors: 8, 8, 8, 8
        1079 => x"08080808",		-- colors: 8, 8, 8, 8
        1080 => x"08080808",		-- colors: 8, 8, 8, 8
        1081 => x"08080808",		-- colors: 8, 8, 8, 8
        1082 => x"08080808",		-- colors: 8, 8, 8, 8
        1083 => x"08080808",		-- colors: 8, 8, 8, 8
        1084 => x"08080808",		-- colors: 8, 8, 8, 8
        1085 => x"08080808",		-- colors: 8, 8, 8, 8
        1086 => x"08080808",		-- colors: 8, 8, 8, 8
        1087 => x"08080808",		-- colors: 8, 8, 8, 8
        1088 => x"08080808",		-- colors: 8, 8, 8, 8
        1089 => x"08080808",		-- colors: 8, 8, 8, 8
        1090 => x"08080808",		-- colors: 8, 8, 8, 8
        1091 => x"08080808",		-- colors: 8, 8, 8, 8
        1092 => x"08080808",		-- colors: 8, 8, 8, 8
        1093 => x"08080808",		-- colors: 8, 8, 8, 8
        1094 => x"08080808",		-- colors: 8, 8, 8, 8
        1095 => x"08080808",		-- colors: 8, 8, 8, 8
        1096 => x"08080808",		-- colors: 8, 8, 8, 8
        1097 => x"08080808",		-- colors: 8, 8, 8, 8
        1098 => x"08080808",		-- colors: 8, 8, 8, 8
        1099 => x"08080808",		-- colors: 8, 8, 8, 8
        1100 => x"08080808",		-- colors: 8, 8, 8, 8
        1101 => x"08080808",		-- colors: 8, 8, 8, 8
        1102 => x"08080808",		-- colors: 8, 8, 8, 8
        1103 => x"08080808",		-- colors: 8, 8, 8, 8
        1104 => x"08080808",		-- colors: 8, 8, 8, 8
        1105 => x"08080808",		-- colors: 8, 8, 8, 8
        1106 => x"08080808",		-- colors: 8, 8, 8, 8
        1107 => x"08080808",		-- colors: 8, 8, 8, 8
        1108 => x"08080808",		-- colors: 8, 8, 8, 8
        1109 => x"08080808",		-- colors: 8, 8, 8, 8
        1110 => x"08080808",		-- colors: 8, 8, 8, 8
        1111 => x"08080808",		-- colors: 8, 8, 8, 8
        1112 => x"08080808",		-- colors: 8, 8, 8, 8
        1113 => x"08080808",		-- colors: 8, 8, 8, 8
        1114 => x"08080808",		-- colors: 8, 8, 8, 8
        1115 => x"08080808",		-- colors: 8, 8, 8, 8
        1116 => x"08080808",		-- colors: 8, 8, 8, 8
        1117 => x"08080808",		-- colors: 8, 8, 8, 8
        1118 => x"08080808",		-- colors: 8, 8, 8, 8
        1119 => x"08080808",		-- colors: 8, 8, 8, 8
        1120 => x"08080808",		-- colors: 8, 8, 8, 8
        1121 => x"08080808",		-- colors: 8, 8, 8, 8
        1122 => x"08080808",		-- colors: 8, 8, 8, 8
        1123 => x"08080808",		-- colors: 8, 8, 8, 8
        1124 => x"08080808",		-- colors: 8, 8, 8, 8
        1125 => x"08080808",		-- colors: 8, 8, 8, 8
        1126 => x"08080808",		-- colors: 8, 8, 8, 8
        1127 => x"08080808",		-- colors: 8, 8, 8, 8

                --  sprite 2
        1128 => x"09090909",		-- colors: 9, 9, 9, 9
        1129 => x"09090909",		-- colors: 9, 9, 9, 9
        1130 => x"09090909",		-- colors: 9, 9, 9, 9
        1131 => x"09090909",		-- colors: 9, 9, 9, 9
        1132 => x"09090909",		-- colors: 9, 9, 9, 9
        1133 => x"09090909",		-- colors: 9, 9, 9, 9
        1134 => x"09090909",		-- colors: 9, 9, 9, 9
        1135 => x"09090909",		-- colors: 9, 9, 9, 9
        1136 => x"09090909",		-- colors: 9, 9, 9, 9
        1137 => x"09090909",		-- colors: 9, 9, 9, 9
        1138 => x"09090909",		-- colors: 9, 9, 9, 9
        1139 => x"09090909",		-- colors: 9, 9, 9, 9
        1140 => x"09090909",		-- colors: 9, 9, 9, 9
        1141 => x"09090909",		-- colors: 9, 9, 9, 9
        1142 => x"09090909",		-- colors: 9, 9, 9, 9
        1143 => x"09090909",		-- colors: 9, 9, 9, 9
        1144 => x"09090909",		-- colors: 9, 9, 9, 9
        1145 => x"09090909",		-- colors: 9, 9, 9, 9
        1146 => x"09090909",		-- colors: 9, 9, 9, 9
        1147 => x"09090909",		-- colors: 9, 9, 9, 9
        1148 => x"09090909",		-- colors: 9, 9, 9, 9
        1149 => x"09090909",		-- colors: 9, 9, 9, 9
        1150 => x"09090909",		-- colors: 9, 9, 9, 9
        1151 => x"09090909",		-- colors: 9, 9, 9, 9
        1152 => x"09090909",		-- colors: 9, 9, 9, 9
        1153 => x"09090909",		-- colors: 9, 9, 9, 9
        1154 => x"09090909",		-- colors: 9, 9, 9, 9
        1155 => x"09090909",		-- colors: 9, 9, 9, 9
        1156 => x"09090909",		-- colors: 9, 9, 9, 9
        1157 => x"09090909",		-- colors: 9, 9, 9, 9
        1158 => x"09090909",		-- colors: 9, 9, 9, 9
        1159 => x"09090909",		-- colors: 9, 9, 9, 9
        1160 => x"09090909",		-- colors: 9, 9, 9, 9
        1161 => x"09090909",		-- colors: 9, 9, 9, 9
        1162 => x"09090909",		-- colors: 9, 9, 9, 9
        1163 => x"09090909",		-- colors: 9, 9, 9, 9
        1164 => x"09090909",		-- colors: 9, 9, 9, 9
        1165 => x"09090909",		-- colors: 9, 9, 9, 9
        1166 => x"09090909",		-- colors: 9, 9, 9, 9
        1167 => x"09090909",		-- colors: 9, 9, 9, 9
        1168 => x"09090909",		-- colors: 9, 9, 9, 9
        1169 => x"09090909",		-- colors: 9, 9, 9, 9
        1170 => x"09090909",		-- colors: 9, 9, 9, 9
        1171 => x"09090909",		-- colors: 9, 9, 9, 9
        1172 => x"09090909",		-- colors: 9, 9, 9, 9
        1173 => x"09090909",		-- colors: 9, 9, 9, 9
        1174 => x"09090909",		-- colors: 9, 9, 9, 9
        1175 => x"09090909",		-- colors: 9, 9, 9, 9
        1176 => x"09090909",		-- colors: 9, 9, 9, 9
        1177 => x"09090909",		-- colors: 9, 9, 9, 9
        1178 => x"09090909",		-- colors: 9, 9, 9, 9
        1179 => x"09090909",		-- colors: 9, 9, 9, 9
        1180 => x"09090909",		-- colors: 9, 9, 9, 9
        1181 => x"09090909",		-- colors: 9, 9, 9, 9
        1182 => x"09090909",		-- colors: 9, 9, 9, 9
        1183 => x"09090909",		-- colors: 9, 9, 9, 9
        1184 => x"09090909",		-- colors: 9, 9, 9, 9
        1185 => x"09090909",		-- colors: 9, 9, 9, 9
        1186 => x"09090909",		-- colors: 9, 9, 9, 9
        1187 => x"09090909",		-- colors: 9, 9, 9, 9
        1188 => x"09090909",		-- colors: 9, 9, 9, 9
        1189 => x"09090909",		-- colors: 9, 9, 9, 9
        1190 => x"09090909",		-- colors: 9, 9, 9, 9
        1191 => x"09090909",		-- colors: 9, 9, 9, 9

                --  sprite 3
        1192 => x"07070707",		-- colors: 7, 7, 7, 7
        1193 => x"07070707",		-- colors: 7, 7, 7, 7
        1194 => x"07070707",		-- colors: 7, 7, 7, 7
        1195 => x"07070707",		-- colors: 7, 7, 7, 7
        1196 => x"07070707",		-- colors: 7, 7, 7, 7
        1197 => x"07070707",		-- colors: 7, 7, 7, 7
        1198 => x"07070707",		-- colors: 7, 7, 7, 7
        1199 => x"07070707",		-- colors: 7, 7, 7, 7
        1200 => x"07070707",		-- colors: 7, 7, 7, 7
        1201 => x"07070707",		-- colors: 7, 7, 7, 7
        1202 => x"07070707",		-- colors: 7, 7, 7, 7
        1203 => x"07070707",		-- colors: 7, 7, 7, 7
        1204 => x"07070707",		-- colors: 7, 7, 7, 7
        1205 => x"07070707",		-- colors: 7, 7, 7, 7
        1206 => x"07070707",		-- colors: 7, 7, 7, 7
        1207 => x"07070707",		-- colors: 7, 7, 7, 7
        1208 => x"07070707",		-- colors: 7, 7, 7, 7
        1209 => x"07070707",		-- colors: 7, 7, 7, 7
        1210 => x"07070707",		-- colors: 7, 7, 7, 7
        1211 => x"07070707",		-- colors: 7, 7, 7, 7
        1212 => x"07070707",		-- colors: 7, 7, 7, 7
        1213 => x"07070707",		-- colors: 7, 7, 7, 7
        1214 => x"07070707",		-- colors: 7, 7, 7, 7
        1215 => x"07070707",		-- colors: 7, 7, 7, 7
        1216 => x"07070707",		-- colors: 7, 7, 7, 7
        1217 => x"07070707",		-- colors: 7, 7, 7, 7
        1218 => x"07070707",		-- colors: 7, 7, 7, 7
        1219 => x"07070707",		-- colors: 7, 7, 7, 7
        1220 => x"0F0F0F0F",		-- colors: 15, 15, 15, 15
        1221 => x"0F0F0F0F",		-- colors: 15, 15, 15, 15
        1222 => x"0F0F0F0F",		-- colors: 15, 15, 15, 15
        1223 => x"0F0F0F0F",		-- colors: 15, 15, 15, 15
        1224 => x"0F0F0F0F",		-- colors: 15, 15, 15, 15
        1225 => x"0F0F0F0F",		-- colors: 15, 15, 15, 15
        1226 => x"0F0F0F0F",		-- colors: 15, 15, 15, 15
        1227 => x"0F0F0F0F",		-- colors: 15, 15, 15, 15
        1228 => x"07070707",		-- colors: 7, 7, 7, 7
        1229 => x"07070707",		-- colors: 7, 7, 7, 7
        1230 => x"07070707",		-- colors: 7, 7, 7, 7
        1231 => x"07070707",		-- colors: 7, 7, 7, 7
        1232 => x"07070707",		-- colors: 7, 7, 7, 7
        1233 => x"07070707",		-- colors: 7, 7, 7, 7
        1234 => x"07070707",		-- colors: 7, 7, 7, 7
        1235 => x"07070707",		-- colors: 7, 7, 7, 7
        1236 => x"07070707",		-- colors: 7, 7, 7, 7
        1237 => x"07070707",		-- colors: 7, 7, 7, 7
        1238 => x"07070707",		-- colors: 7, 7, 7, 7
        1239 => x"07070707",		-- colors: 7, 7, 7, 7
        1240 => x"07070707",		-- colors: 7, 7, 7, 7
        1241 => x"07070707",		-- colors: 7, 7, 7, 7
        1242 => x"07070707",		-- colors: 7, 7, 7, 7
        1243 => x"07070707",		-- colors: 7, 7, 7, 7
        1244 => x"07070707",		-- colors: 7, 7, 7, 7
        1245 => x"07070707",		-- colors: 7, 7, 7, 7
        1246 => x"07070707",		-- colors: 7, 7, 7, 7
        1247 => x"07070707",		-- colors: 7, 7, 7, 7
        1248 => x"07070707",		-- colors: 7, 7, 7, 7
        1249 => x"07070707",		-- colors: 7, 7, 7, 7
        1250 => x"07070707",		-- colors: 7, 7, 7, 7
        1251 => x"07070707",		-- colors: 7, 7, 7, 7
        1252 => x"07070707",		-- colors: 7, 7, 7, 7
        1253 => x"07070707",		-- colors: 7, 7, 7, 7
        1254 => x"07070707",		-- colors: 7, 7, 7, 7
        1255 => x"07070707",		-- colors: 7, 7, 7, 7

                --  sprite 4
        1256 => x"08080808",		-- colors: 8, 8, 8, 8
        1257 => x"08080A0B",		-- colors: 8, 8, 10, 11
        1258 => x"0A080808",		-- colors: 10, 8, 8, 8
        1259 => x"08080808",		-- colors: 8, 8, 8, 8
        1260 => x"08080C0A",		-- colors: 8, 8, 12, 10
        1261 => x"0A0A0A0A",		-- colors: 10, 10, 10, 10
        1262 => x"0A0A0A0A",		-- colors: 10, 10, 10, 10
        1263 => x"08080808",		-- colors: 8, 8, 8, 8
        1264 => x"080D0A0A",		-- colors: 8, 13, 10, 10
        1265 => x"0A0A0A0A",		-- colors: 10, 10, 10, 10
        1266 => x"0A0A0A0A",		-- colors: 10, 10, 10, 10
        1267 => x"0A080808",		-- colors: 10, 8, 8, 8
        1268 => x"080D0A0A",		-- colors: 8, 13, 10, 10
        1269 => x"0A0A0A0A",		-- colors: 10, 10, 10, 10
        1270 => x"0A0A0A0A",		-- colors: 10, 10, 10, 10
        1271 => x"0A0A0808",		-- colors: 10, 10, 8, 8
        1272 => x"08080D0A",		-- colors: 8, 8, 13, 10
        1273 => x"0A0A0A0A",		-- colors: 10, 10, 10, 10
        1274 => x"0A0A0A0A",		-- colors: 10, 10, 10, 10
        1275 => x"0A0A0A08",		-- colors: 10, 10, 10, 8
        1276 => x"0E0D0A0A",		-- colors: 14, 13, 10, 10
        1277 => x"0A0A0A0A",		-- colors: 10, 10, 10, 10
        1278 => x"0A0A0A0A",		-- colors: 10, 10, 10, 10
        1279 => x"0A0A0A08",		-- colors: 10, 10, 10, 8
        1280 => x"0D0A0A0A",		-- colors: 13, 10, 10, 10
        1281 => x"0A0A0A0A",		-- colors: 10, 10, 10, 10
        1282 => x"0A0A0A0A",		-- colors: 10, 10, 10, 10
        1283 => x"0A0A0808",		-- colors: 10, 10, 8, 8
        1284 => x"0D0A0A0A",		-- colors: 13, 10, 10, 10
        1285 => x"0A0A0A0A",		-- colors: 10, 10, 10, 10
        1286 => x"0A0A0A0A",		-- colors: 10, 10, 10, 10
        1287 => x"0A0A0808",		-- colors: 10, 10, 8, 8
        1288 => x"0D0A0A0A",		-- colors: 13, 10, 10, 10
        1289 => x"0A0A0A0A",		-- colors: 10, 10, 10, 10
        1290 => x"0A0A0A0A",		-- colors: 10, 10, 10, 10
        1291 => x"0A0A0808",		-- colors: 10, 10, 8, 8
        1292 => x"080D0A0A",		-- colors: 8, 13, 10, 10
        1293 => x"0A0A0A0A",		-- colors: 10, 10, 10, 10
        1294 => x"0A0A0A0A",		-- colors: 10, 10, 10, 10
        1295 => x"0A0A0808",		-- colors: 10, 10, 8, 8
        1296 => x"080D0A0A",		-- colors: 8, 13, 10, 10
        1297 => x"0A0A0A0A",		-- colors: 10, 10, 10, 10
        1298 => x"0A0A0A0A",		-- colors: 10, 10, 10, 10
        1299 => x"08080808",		-- colors: 8, 8, 8, 8
        1300 => x"080D0A0A",		-- colors: 8, 13, 10, 10
        1301 => x"0A0A0A0A",		-- colors: 10, 10, 10, 10
        1302 => x"0A0A0A08",		-- colors: 10, 10, 10, 8
        1303 => x"08080808",		-- colors: 8, 8, 8, 8
        1304 => x"080D0A0A",		-- colors: 8, 13, 10, 10
        1305 => x"0A0A0A0A",		-- colors: 10, 10, 10, 10
        1306 => x"0A0A0A08",		-- colors: 10, 10, 10, 8
        1307 => x"08080808",		-- colors: 8, 8, 8, 8
        1308 => x"080E0D0A",		-- colors: 8, 14, 13, 10
        1309 => x"0D0D0A0A",		-- colors: 13, 13, 10, 10
        1310 => x"0A0A0808",		-- colors: 10, 10, 8, 8
        1311 => x"08080808",		-- colors: 8, 8, 8, 8
        1312 => x"0808080E",		-- colors: 8, 8, 8, 14
        1313 => x"08080A0A",		-- colors: 8, 8, 10, 10
        1314 => x"0A080808",		-- colors: 10, 8, 8, 8
        1315 => x"08080808",		-- colors: 8, 8, 8, 8
        1316 => x"08080808",		-- colors: 8, 8, 8, 8
        1317 => x"08080808",		-- colors: 8, 8, 8, 8
        1318 => x"08080808",		-- colors: 8, 8, 8, 8
        1319 => x"08080808",		-- colors: 8, 8, 8, 8

others => x"00000000"
	);


begin

	process(i_clk)
	begin
		if rising_edge(i_clk) then
			-- memory write --
			if i_we = '1' then
				mem(to_integer(unsigned(i_w_addr))) <= i_data;
			end if;
			-- memory read -- 
			o_data <= mem(to_integer(unsigned(i_r_addr)));
			
		end if; 
	end process;

end architecture arch;
